module dpram_2048x20
(
  // Clock & reset
  input         reset,
  input         clock,
  // Port A : micro-instruction fetch
  input         rden_a,
  input  [10:0] address_a,
  output [19:0] q_a,
  // Port B : m68k registers read/write
  input   [1:0] wren_b,
  input  [10:0] address_b,
  input  [15:0] data_b,
  output [15:0] q_b
);

// Inferred block ROM and RAM
reg  [15:0] r_mem_blk [0:2047];

reg  [19:0] r_q_a;
reg  [15:0] r_q_b;

// Port A (read only)
always@(posedge reset or posedge clock) begin
  if (reset)
    r_q_a <= 20'hC0458; // NOP instruction
  else if (rden_a) begin
    case(address_a)
      11'h000 : r_q_a <= 20'b11000000010001011000; // C0458 NOP
      11'h001 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h002 : r_q_a <= 20'b00000000000000000100; // 00004 LOOP #16
      11'h003 : r_q_a <= 20'b10100000010101000111; // A0547 WRW RH[CNT]
      11'h004 : r_q_a <= 20'b10100000010001000111; // A0447 WRW RL[CNT]
      11'h005 : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h006 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h007 : r_q_a <= 20'b10000011010001000110; // 83446 STW VECL
      11'h008 : r_q_a <= 20'b10000101010110000111; // 85587 LDW (VEC)+
      11'h009 : r_q_a <= 20'b10100000010101001111; // A054F WRW SSPH
      11'h00A : r_q_a <= 20'b10100011010101000011; // A3543 STW A7H
      11'h00B : r_q_a <= 20'b10000101010110000111; // 85587 LDW (VEC)+
      11'h00C : r_q_a <= 20'b10100000010001001111; // A044F WRW SSPL
      11'h00D : r_q_a <= 20'b10100011010001000011; // A3443 STW A7L
      11'h00E : r_q_a <= 20'b01000010011100000100; // 42704 LIT #2704
      11'h00F : r_q_a <= 20'b00101110011011010000; // 2E6D0 CALL Resume_Exec
      11'h010 : r_q_a <= 20'b10000000010110000010; // 80582 FTI (PC)+
      11'h011 : r_q_a <= 20'b10000101010010001100; // 8548C LDW DECJ
      11'h012 : r_q_a <= 20'b00101111000000000000; // 2F000 CALL 0000(T)
      11'h013 : r_q_a <= 20'b00111011100000010000; // 3B810 JUMPN I_SR,Decode
      11'h014 : r_q_a <= 20'b00111101000000011111; // 3D01F JUMP T_SR,Trap_Trace
      11'h015 : r_q_a <= 20'b00110000000000100010; // 30022 JUMP A_SR,Trap_Address
      11'h016 : r_q_a <= 20'b00101110011010111110; // 2E6BE CALL Enter_Super
      11'h017 : r_q_a <= 20'b00101110011010100001; // 2E6A1 CALL PC_SR_to_Stack
      11'h018 : r_q_a <= 20'b00101110011011001011; // 2E6CB CALL SR_Super
      11'h019 : r_q_a <= 20'b01000010000011111111; // 420FF LIT #20FF
      11'h01A : r_q_a <= 20'b11000011010001001010; // C344A ANDW
      11'h01B : r_q_a <= 20'b10000101010010000110; // 85486 LDW VECL
      11'h01C : r_q_a <= 20'b11000011010001011010; // C345A ORW
      11'h01D : r_q_a <= 20'b00101110011011010000; // 2E6D0 CALL Resume_Exec
      11'h01E : r_q_a <= 20'b00111110000000010000; // 3E010 JUMP Decode
      11'h01F : r_q_a <= 20'b01000000000000100100; // 40024 LIT #0024
      11'h020 : r_q_a <= 20'b00101110000001000001; // 2E041 CALL Trap_Processing
      11'h021 : r_q_a <= 20'b00111110000000010000; // 3E010 JUMP Decode
      11'h022 : r_q_a <= 20'b01000000000000001100; // 4000C LIT #000C
      11'h023 : r_q_a <= 20'b10000011010001000110; // 83446 STW VECL
      11'h024 : r_q_a <= 20'b00101110011010111110; // 2E6BE CALL Enter_Super
      11'h025 : r_q_a <= 20'b00101110011010100001; // 2E6A1 CALL PC_SR_to_Stack
      11'h026 : r_q_a <= 20'b10000101010010000111; // 85487 LDW CPUS
      11'h027 : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h028 : r_q_a <= 20'b10000101010010000111; // 85487 LDW CPUS
      11'h029 : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h02A : r_q_a <= 20'b10000101010010000111; // 85487 LDW CPUS
      11'h02B : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h02C : r_q_a <= 20'b10000101010010000111; // 85487 LDW CPUS
      11'h02D : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h02E : r_q_a <= 20'b00101110011010101110; // 2E6AE CALL EA2_to_SP
      11'h02F : r_q_a <= 20'b00101110011011001011; // 2E6CB CALL SR_Super
      11'h030 : r_q_a <= 20'b00101110011011010000; // 2E6D0 CALL Resume_Exec
      11'h031 : r_q_a <= 20'b00111110000000010000; // 3E010 JUMP Decode
      11'h032 : r_q_a <= 20'b01000000000000101100; // 4002C LIT #002C
      11'h033 : r_q_a <= 20'b00111110000001000001; // 3E041 JUMP Trap_Processing
      11'h034 : r_q_a <= 20'b01000000000000101000; // 40028 LIT #0028
      11'h035 : r_q_a <= 20'b00111110000001000001; // 3E041 JUMP Trap_Processing
      11'h036 : r_q_a <= 20'b01000000000000010100; // 40014 LIT #0014
      11'h037 : r_q_a <= 20'b00111110000001000001; // 3E041 JUMP Trap_Processing
      11'h038 : r_q_a <= 20'b01000000000000100000; // 40020 LIT #0020
      11'h039 : r_q_a <= 20'b00111110000000111011; // 3E03B JUMP Trap_Processing2
      11'h03A : r_q_a <= 20'b01000000000000010000; // 40010 LIT #0010
      11'h03B : r_q_a <= 20'b10000101010010000101; // 85485 LDW PCH
      11'h03C : r_q_a <= 20'b10000101010010000100; // 85484 LDW PCL
      11'h03D : r_q_a <= 20'b01001111111111111110; // 4FFFE LIT #FFFE
      11'h03E : r_q_a <= 20'b00101110011010010000; // 2E690 CALL AddVal
      11'h03F : r_q_a <= 20'b10000011010001000101; // 83445 STW PCH
      11'h040 : r_q_a <= 20'b10000011010001000100; // 83444 STW PCL
      11'h041 : r_q_a <= 20'b10000011010001000110; // 83446 STW VECL
      11'h042 : r_q_a <= 20'b00101110011010111110; // 2E6BE CALL Enter_Super
      11'h043 : r_q_a <= 20'b00101110011010100001; // 2E6A1 CALL PC_SR_to_Stack
      11'h044 : r_q_a <= 20'b00101110011011001011; // 2E6CB CALL SR_Super
      11'h045 : r_q_a <= 20'b00111110011011010000; // 3E6D0 JUMP Resume_Exec
      11'h046 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h047 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h048 : r_q_a <= 20'b11000011001001011010; // C325A ORB.
      11'h049 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h04A : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h04B : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h04C : r_q_a <= 20'b10000101000010001111; // 8508F LDB SR
      11'h04D : r_q_a <= 20'b11000011000001011010; // C305A ORB
      11'h04E : r_q_a <= 20'b10010011000001001111; // 9304F STB SR; RTS
      11'h04F : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h050 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h051 : r_q_a <= 20'b11000011011001011010; // C365A ORW.
      11'h052 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h053 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h054 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h055 : r_q_a <= 20'b10000101010010001111; // 8548F LDW SR
      11'h056 : r_q_a <= 20'b11000011010001011010; // C345A ORW
      11'h057 : r_q_a <= 20'b10000011010001001111; // 8344F STW SR
      11'h058 : r_q_a <= 20'b00111110011011001000; // 3E6C8 JUMP Leave_Super
      11'h059 : r_q_a <= 20'b00101110011000101010; // 2E62A CALL EA1_RL_to_TMP1
      11'h05A : r_q_a <= 20'b11000011011001011010; // C365A ORW.
      11'h05B : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h05C : r_q_a <= 20'b10100101010110001100; // A558C LDW TMP1H
      11'h05D : r_q_a <= 20'b11000011101001011010; // C3A5A ORL.
      11'h05E : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h05F : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h060 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h061 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h062 : r_q_a <= 20'b11000011001001001010; // C324A ANDB.
      11'h063 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h064 : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h065 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h066 : r_q_a <= 20'b10000101000010001111; // 8508F LDB SR
      11'h067 : r_q_a <= 20'b11000011000001001010; // C304A ANDB
      11'h068 : r_q_a <= 20'b10010011000001001111; // 9304F STB SR; RTS
      11'h069 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h06A : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h06B : r_q_a <= 20'b11000011011001001010; // C364A ANDW.
      11'h06C : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h06D : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h06E : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h06F : r_q_a <= 20'b10000101010010001111; // 8548F LDW SR
      11'h070 : r_q_a <= 20'b11000011010001001010; // C344A ANDW
      11'h071 : r_q_a <= 20'b10000011010001001111; // 8344F STW SR
      11'h072 : r_q_a <= 20'b00111110011011001000; // 3E6C8 JUMP Leave_Super
      11'h073 : r_q_a <= 20'b00101110011000101010; // 2E62A CALL EA1_RL_to_TMP1
      11'h074 : r_q_a <= 20'b11000011011001001010; // C364A ANDW.
      11'h075 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h076 : r_q_a <= 20'b10100101010110001100; // A558C LDW TMP1H
      11'h077 : r_q_a <= 20'b11000011101001001010; // C3A4A ANDL.
      11'h078 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h079 : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h07A : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h07B : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h07C : r_q_a <= 20'b11000011001000101011; // C322B SUBB.
      11'h07D : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h07E : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h07F : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h080 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h081 : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h082 : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h083 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h084 : r_q_a <= 20'b00101110011000101010; // 2E62A CALL EA1_RL_to_TMP1
      11'h085 : r_q_a <= 20'b11000011011000101110; // C362E SUBW.
      11'h086 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h087 : r_q_a <= 20'b10100101010110001100; // A558C LDW TMP1H
      11'h088 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h089 : r_q_a <= 20'b11000011101000111110; // C3A3E SUBCL.
      11'h08A : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h08B : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h08C : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h08D : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h08E : r_q_a <= 20'b11000011001000001010; // C320A ADDB.
      11'h08F : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h090 : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h091 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h092 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h093 : r_q_a <= 20'b11000011011000001010; // C360A ADDW.
      11'h094 : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h095 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h096 : r_q_a <= 20'b00101110011000101010; // 2E62A CALL EA1_RL_to_TMP1
      11'h097 : r_q_a <= 20'b11000011011000001010; // C360A ADDW.
      11'h098 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h099 : r_q_a <= 20'b10100101010110001100; // A558C LDW TMP1H
      11'h09A : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h09B : r_q_a <= 20'b11000011101000011010; // C3A1A ADDCL.
      11'h09C : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h09D : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h09E : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h09F : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h0A0 : r_q_a <= 20'b11000011001101001010; // C334A BANDB.
      11'h0A1 : r_q_a <= 20'b01100000100000010000; // 60810 FLAG --*--,CIN=CLR
      11'h0A2 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h0A3 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h0A4 : r_q_a <= 20'b11000101010001010010; // C5452 OVER
      11'h0A5 : r_q_a <= 20'b11000101010001010010; // C5452 OVER
      11'h0A6 : r_q_a <= 20'b11000011001101001010; // C334A BANDB.
      11'h0A7 : r_q_a <= 20'b01100000100000010000; // 60810 FLAG --*--,CIN=CLR
      11'h0A8 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h0A9 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h0AA : r_q_a <= 20'b11000101010001011000; // C5458 DUP
      11'h0AB : r_q_a <= 20'b10100101010010000010; // A5482 LDW RL[EA1]
      11'h0AC : r_q_a <= 20'b11000011011101001010; // C374A BANDW.
      11'h0AD : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h0AE : r_q_a <= 20'b10100101010110000010; // A5582 LDW RH[EA1]
      11'h0AF : r_q_a <= 20'b11000011101101001010; // C3B4A BANDL.
      11'h0B0 : r_q_a <= 20'b01100000100000010000; // 60810 FLAG --*--,CIN=CLR
      11'h0B1 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h0B2 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h0B3 : r_q_a <= 20'b00101110000010100011; // 2E0A3 CALL Op_BTSTB_call
      11'h0B4 : r_q_a <= 20'b11000011000101101010; // C316A BXORB
      11'h0B5 : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h0B6 : r_q_a <= 20'b00101110000010101001; // 2E0A9 CALL Op_BTSTL_i
      11'h0B7 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h0B8 : r_q_a <= 20'b11000101010001011000; // C5458 DUP
      11'h0B9 : r_q_a <= 20'b10100101010010000010; // A5482 LDW RL[EA1]
      11'h0BA : r_q_a <= 20'b11000011010101101010; // C356A BXORW
      11'h0BB : r_q_a <= 20'b10100011010001000010; // A3442 STW RL[EA1]
      11'h0BC : r_q_a <= 20'b10100101010110000010; // A5582 LDW RH[EA1]
      11'h0BD : r_q_a <= 20'b11000011100101101010; // C396A BXORL
      11'h0BE : r_q_a <= 20'b10110011010101000010; // B3542 STW RH[EA1]; RTS
      11'h0BF : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h0C0 : r_q_a <= 20'b00101110000010100011; // 2E0A3 CALL Op_BTSTB_call
      11'h0C1 : r_q_a <= 20'b11000011000101001011; // C314B BMSKB
      11'h0C2 : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h0C3 : r_q_a <= 20'b00101110000010101001; // 2E0A9 CALL Op_BTSTL_i
      11'h0C4 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h0C5 : r_q_a <= 20'b11000101010001011000; // C5458 DUP
      11'h0C6 : r_q_a <= 20'b10100101010010000010; // A5482 LDW RL[EA1]
      11'h0C7 : r_q_a <= 20'b11000011010101001011; // C354B BMSKW
      11'h0C8 : r_q_a <= 20'b10100011010001000010; // A3442 STW RL[EA1]
      11'h0C9 : r_q_a <= 20'b10100101010110000010; // A5582 LDW RH[EA1]
      11'h0CA : r_q_a <= 20'b11000011100101001011; // C394B BMSKL
      11'h0CB : r_q_a <= 20'b10110011010101000010; // B3542 STW RH[EA1]; RTS
      11'h0CC : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h0CD : r_q_a <= 20'b00101110000010100011; // 2E0A3 CALL Op_BTSTB_call
      11'h0CE : r_q_a <= 20'b11000011000101011010; // C315A BORB
      11'h0CF : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h0D0 : r_q_a <= 20'b00101110000010101001; // 2E0A9 CALL Op_BTSTL_i
      11'h0D1 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h0D2 : r_q_a <= 20'b11000101010001011000; // C5458 DUP
      11'h0D3 : r_q_a <= 20'b10100101010010000010; // A5482 LDW RL[EA1]
      11'h0D4 : r_q_a <= 20'b11000011010101011010; // C355A BORW
      11'h0D5 : r_q_a <= 20'b10100011010001000010; // A3442 STW RL[EA1]
      11'h0D6 : r_q_a <= 20'b10100101010110000010; // A5582 LDW RH[EA1]
      11'h0D7 : r_q_a <= 20'b11000011100101011010; // C395A BORL
      11'h0D8 : r_q_a <= 20'b10110011010101000010; // B3542 STW RH[EA1]; RTS
      11'h0D9 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h0DA : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h0DB : r_q_a <= 20'b11000011001001101010; // C326A XORB.
      11'h0DC : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h0DD : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h0DE : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h0DF : r_q_a <= 20'b10000101000010001111; // 8508F LDB SR
      11'h0E0 : r_q_a <= 20'b11000011000001101010; // C306A XORB
      11'h0E1 : r_q_a <= 20'b10010011000001001111; // 9304F STB SR; RTS
      11'h0E2 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h0E3 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h0E4 : r_q_a <= 20'b11000011011001101010; // C366A XORW.
      11'h0E5 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h0E6 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h0E7 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h0E8 : r_q_a <= 20'b10000101010010001111; // 8548F LDW SR
      11'h0E9 : r_q_a <= 20'b11000011010001101010; // C346A XORW
      11'h0EA : r_q_a <= 20'b10000011010001001111; // 8344F STW SR
      11'h0EB : r_q_a <= 20'b00111110011011001000; // 3E6C8 JUMP Leave_Super
      11'h0EC : r_q_a <= 20'b00101110011000101010; // 2E62A CALL EA1_RL_to_TMP1
      11'h0ED : r_q_a <= 20'b11000011011001101010; // C366A XORW.
      11'h0EE : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h0EF : r_q_a <= 20'b10100101010110001100; // A558C LDW TMP1H
      11'h0F0 : r_q_a <= 20'b11000011101001101010; // C3A6A XORL.
      11'h0F1 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h0F2 : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h0F3 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h0F4 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h0F5 : r_q_a <= 20'b11000011001000101011; // C322B SUBB.
      11'h0F6 : r_q_a <= 20'b01100000100010010101; // 60895 FLAG -****,CIN=CLR
      11'h0F7 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h0F8 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h0F9 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h0FA : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h0FB : r_q_a <= 20'b01100000100010010101; // 60895 FLAG -****,CIN=CLR
      11'h0FC : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h0FD : r_q_a <= 20'b00101110011000101010; // 2E62A CALL EA1_RL_to_TMP1
      11'h0FE : r_q_a <= 20'b11000011011000101110; // C362E SUBW.
      11'h0FF : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h100 : r_q_a <= 20'b10100101010110001100; // A558C LDW TMP1H
      11'h101 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h102 : r_q_a <= 20'b11000011101000111110; // C3A3E SUBCL.
      11'h103 : r_q_a <= 20'b01100000100010010101; // 60895 FLAG -****,CIN=CLR
      11'h104 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h105 : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h106 : r_q_a <= 20'b00111110000010011111; // 3E09F JUMP Op_BTSTB_jmp
      11'h107 : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h108 : r_q_a <= 20'b00111110000010101010; // 3E0AA JUMP Op_BTSTL_jmp
      11'h109 : r_q_a <= 20'b00101110011011100010; // 2E6E2 CALL Calc_d16_An_EA1
      11'h10A : r_q_a <= 20'b00111110000100010110; // 3E116 JUMP Op_MOVEPW_r_jmp
      11'h10B : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h10C : r_q_a <= 20'b00111110000010110011; // 3E0B3 JUMP Op_BCHGB_jmp
      11'h10D : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h10E : r_q_a <= 20'b11000101010001011000; // C5458 DUP
      11'h10F : r_q_a <= 20'b00101110000010101010; // 2E0AA CALL Op_BTSTL_jmp
      11'h110 : r_q_a <= 20'b00111110000010111000; // 3E0B8 JUMP Op_BCHGL_jmp
      11'h111 : r_q_a <= 20'b00101110011011100010; // 2E6E2 CALL Calc_d16_An_EA1
      11'h112 : r_q_a <= 20'b10000101110110000100; // 85D84 LDH (EA1)+
      11'h113 : r_q_a <= 20'b10000101100110000100; // 85984 LDL (EA1)+
      11'h114 : r_q_a <= 20'b11000011010001011010; // C345A ORW
      11'h115 : r_q_a <= 20'b10100011010101000100; // A3544 STW DH[EA2]
      11'h116 : r_q_a <= 20'b10000101110110000100; // 85D84 LDH (EA1)+
      11'h117 : r_q_a <= 20'b10000101100110000000; // 85980 LDL (EA1)
      11'h118 : r_q_a <= 20'b11000011010001011010; // C345A ORW
      11'h119 : r_q_a <= 20'b10110011010001000100; // B3444 STW DL[EA2]; RTS
      11'h11A : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h11B : r_q_a <= 20'b00111110000011000000; // 3E0C0 JUMP Op_BCLRB_jmp
      11'h11C : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h11D : r_q_a <= 20'b11000101010001011000; // C5458 DUP
      11'h11E : r_q_a <= 20'b00101110000010101010; // 2E0AA CALL Op_BTSTL_jmp
      11'h11F : r_q_a <= 20'b00111110000011000101; // 3E0C5 JUMP Op_BCLRL_jmp
      11'h120 : r_q_a <= 20'b00101110011011100010; // 2E6E2 CALL Calc_d16_An_EA1
      11'h121 : r_q_a <= 20'b00111110000100101101; // 3E12D JUMP Op_MOVEPW_m_jmp
      11'h122 : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h123 : r_q_a <= 20'b00111110000011001101; // 3E0CD JUMP Op_BSETB_jmp
      11'h124 : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h125 : r_q_a <= 20'b11000101010001011000; // C5458 DUP
      11'h126 : r_q_a <= 20'b00101110000010101010; // 2E0AA CALL Op_BTSTL_jmp
      11'h127 : r_q_a <= 20'b00111110000011010010; // 3E0D2 JUMP Op_BSETL_jmp
      11'h128 : r_q_a <= 20'b00101110011011100010; // 2E6E2 CALL Calc_d16_An_EA1
      11'h129 : r_q_a <= 20'b10100101010110000100; // A5584 LDW DH[EA2]
      11'h12A : r_q_a <= 20'b11000101010001011000; // C5458 DUP
      11'h12B : r_q_a <= 20'b10000011110101000100; // 83D44 STH (EA1)+
      11'h12C : r_q_a <= 20'b10000011100101000100; // 83944 STL (EA1)+
      11'h12D : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h12E : r_q_a <= 20'b11000101010001011000; // C5458 DUP
      11'h12F : r_q_a <= 20'b10000011110101000100; // 83D44 STH (EA1)+
      11'h130 : r_q_a <= 20'b10010011100101000000; // 93940 STL (EA1); RTS
      11'h131 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h132 : r_q_a <= 20'b11000000001001011000; // C0258 TSTB.
      11'h133 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h134 : r_q_a <= 20'b00111110011001101010; // 3E66A JUMP EA2_Write_B
      11'h135 : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h136 : r_q_a <= 20'b11000000011001011000; // C0658 TSTW.
      11'h137 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h138 : r_q_a <= 20'b11000000101001011000; // C0A58 TSTL.
      11'h139 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h13A : r_q_a <= 20'b00111110011010000000; // 3E680 JUMP EA2_Write_L
      11'h13B : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h13C : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h13D : r_q_a <= 20'b00111110011010000000; // 3E680 JUMP EA2_Write_L
      11'h13E : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h13F : r_q_a <= 20'b11000000011001011000; // C0658 TSTW.
      11'h140 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h141 : r_q_a <= 20'b00111110011001110011; // 3E673 JUMP EA2_Write_W
      11'h142 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h143 : r_q_a <= 20'b00111110011001110011; // 3E673 JUMP EA2_Write_W
      11'h144 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h145 : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h146 : r_q_a <= 20'b11000000001000111100; // C023C NEGCB.
      11'h147 : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h148 : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h149 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h14A : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h14B : r_q_a <= 20'b11000000011000111100; // C063C NEGCW.
      11'h14C : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h14D : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h14E : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h14F : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h150 : r_q_a <= 20'b11000000011000111100; // C063C NEGCW.
      11'h151 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h152 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h153 : r_q_a <= 20'b11000000101000111100; // C0A3C NEGCL.
      11'h154 : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h155 : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h156 : r_q_a <= 20'b10000101010010001111; // 8548F LDW SR
      11'h157 : r_q_a <= 20'b00111110011001000110; // 3E646 JUMP EA1_Write_W
      11'h158 : r_q_a <= 20'b01100000000100111010; // 6013A FLAG -0100,CIN=KEEP
      11'h159 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h15A : r_q_a <= 20'b00111110011000111101; // 3E63D JUMP EA1_Write_B
      11'h15B : r_q_a <= 20'b01100000000100111010; // 6013A FLAG -0100,CIN=KEEP
      11'h15C : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h15D : r_q_a <= 20'b00111110011001000110; // 3E646 JUMP EA1_Write_W
      11'h15E : r_q_a <= 20'b01100000000100111010; // 6013A FLAG -0100,CIN=KEEP
      11'h15F : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h160 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h161 : r_q_a <= 20'b00111110011001001111; // 3E64F JUMP EA1_Write_L
      11'h162 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h163 : r_q_a <= 20'b11000000001000101100; // C022C NEGB.
      11'h164 : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h165 : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h166 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h167 : r_q_a <= 20'b11000000011000101100; // C062C NEGW.
      11'h168 : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h169 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h16A : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h16B : r_q_a <= 20'b11000000011000101100; // C062C NEGW.
      11'h16C : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h16D : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h16E : r_q_a <= 20'b11000000101000111100; // C0A3C NEGCL.
      11'h16F : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h170 : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h171 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h172 : r_q_a <= 20'b10010011000001001111; // 9304F STB SR; RTS
      11'h173 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h174 : r_q_a <= 20'b11000000001001111010; // C027A NOTB.
      11'h175 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h176 : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h177 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h178 : r_q_a <= 20'b11000000011001111010; // C067A NOTW.
      11'h179 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h17A : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h17B : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h17C : r_q_a <= 20'b11000000011001111010; // C067A NOTW.
      11'h17D : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h17E : r_q_a <= 20'b11000000101001111010; // C0A7A NOTL.
      11'h17F : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h180 : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h181 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h182 : r_q_a <= 20'b10000011010001001111; // 8344F STW SR
      11'h183 : r_q_a <= 20'b00111110011011001000; // 3E6C8 JUMP Leave_Super
      11'h184 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h185 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h186 : r_q_a <= 20'b00101110001011001101; // 2E2CD CALL SBCD_Calc
      11'h187 : r_q_a <= 20'b01100000100011010000; // 608D0 FLAG -*#--,CIN=CLR
      11'h188 : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h189 : r_q_a <= 20'b00101110011000110000; // 2E630 CALL EA1_Calc
      11'h18A : r_q_a <= 20'b00101110011010110010; // 2E6B2 CALL SP_to_EA2
      11'h18B : r_q_a <= 20'b10000101010010000000; // 85480 LDW EA1L
      11'h18C : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h18D : r_q_a <= 20'b10000101010010000001; // 85481 LDW EA1H
      11'h18E : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h18F : r_q_a <= 20'b00111110011010101110; // 3E6AE JUMP EA2_to_SP
      11'h190 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h191 : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h192 : r_q_a <= 20'b01100000100000001010; // 6080A FLAG ---00,CIN=CLR
      11'h193 : r_q_a <= 20'b11000000011001011000; // C0658 TSTW.
      11'h194 : r_q_a <= 20'b10100011010001000000; // A3440 STW DL[EA1]
      11'h195 : r_q_a <= 20'b11000000101001011000; // C0A58 TSTL.
      11'h196 : r_q_a <= 20'b01100000100010010000; // 60890 FLAG -**--,CIN=CLR
      11'h197 : r_q_a <= 20'b10110011010101000000; // B3540 STW DH[EA1]; RTS
      11'h198 : r_q_a <= 20'b11000000011001011000; // C0658 TSTW.
      11'h199 : r_q_a <= 20'b01100000100010010000; // 60890 FLAG -**--,CIN=CLR
      11'h19A : r_q_a <= 20'b10110011010001000000; // B3440 STW DL[EA1]; RTS
      11'h19B : r_q_a <= 20'b11000000001001011000; // C0258 TSTB.
      11'h19C : r_q_a <= 20'b01100000100010010000; // 60890 FLAG -**--,CIN=CLR
      11'h19D : r_q_a <= 20'b10110011000001000000; // B3040 STB DL[EA1]; RTS
      11'h19E : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h19F : r_q_a <= 20'b00101110011000110000; // 2E630 CALL EA1_Calc
      11'h1A0 : r_q_a <= 20'b00000000000110100100; // 001A4 LOOP #16
      11'h1A1 : r_q_a <= 20'b00110100100110100100; // 349A4 JUMPN T[0],NoMoveW_m
      11'h1A2 : r_q_a <= 20'b10100101010010000111; // A5487 LDW RL[CNT]
      11'h1A3 : r_q_a <= 20'b10000011010101000100; // 83544 STW (EA1)+
      11'h1A4 : r_q_a <= 20'b11000100010011000000; // C44C0 RSHW
      11'h1A5 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h1A6 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h1A7 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h1A8 : r_q_a <= 20'b00000000000110101100; // 001AC LOOP #16
      11'h1A9 : r_q_a <= 20'b00110100100110101100; // 349AC JUMPN T[0],NoMoveW_mpd
      11'h1AA : r_q_a <= 20'b10100101010010000111; // A5487 LDW RL[CNT]
      11'h1AB : r_q_a <= 20'b10000011010101001000; // 83548 STW -(EA1)
      11'h1AC : r_q_a <= 20'b11000100010011000000; // C44C0 RSHW
      11'h1AD : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h1AE : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h1AF : r_q_a <= 20'b01001111111100000000; // 4FF00 LIT #FF00
      11'h1B0 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h1B1 : r_q_a <= 20'b11000000001001011000; // C0258 TSTB.
      11'h1B2 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h1B3 : r_q_a <= 20'b00111001000110110110; // 391B6 JUMP N_SR,Op_EXTW_Neg
      11'h1B4 : r_q_a <= 20'b11000011010001001011; // C344B MSKW
      11'h1B5 : r_q_a <= 20'b10110011010001000000; // B3440 STW DL[EA1]; RTS
      11'h1B6 : r_q_a <= 20'b11000011010001011010; // C345A ORW
      11'h1B7 : r_q_a <= 20'b10110011010001000000; // B3440 STW DL[EA1]; RTS
      11'h1B8 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h1B9 : r_q_a <= 20'b00101110011000110000; // 2E630 CALL EA1_Calc
      11'h1BA : r_q_a <= 20'b00000000000111000000; // 001C0 LOOP #16
      11'h1BB : r_q_a <= 20'b00110100100111000000; // 349C0 JUMPN T[0],NoMoveL_m
      11'h1BC : r_q_a <= 20'b10100101010110000111; // A5587 LDW RH[CNT]
      11'h1BD : r_q_a <= 20'b10000011010101000100; // 83544 STW (EA1)+
      11'h1BE : r_q_a <= 20'b10100101010010000111; // A5487 LDW RL[CNT]
      11'h1BF : r_q_a <= 20'b10000011010101000100; // 83544 STW (EA1)+
      11'h1C0 : r_q_a <= 20'b11000100010011000000; // C44C0 RSHW
      11'h1C1 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h1C2 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h1C3 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h1C4 : r_q_a <= 20'b00000000000111001010; // 001CA LOOP #16
      11'h1C5 : r_q_a <= 20'b00110100100111001010; // 349CA JUMPN T[0],NoMoveL_mpd
      11'h1C6 : r_q_a <= 20'b10100101010010000111; // A5487 LDW RL[CNT]
      11'h1C7 : r_q_a <= 20'b10000011010101001000; // 83548 STW -(EA1)
      11'h1C8 : r_q_a <= 20'b10100101010110000111; // A5587 LDW RH[CNT]
      11'h1C9 : r_q_a <= 20'b10000011010101001000; // 83548 STW -(EA1)
      11'h1CA : r_q_a <= 20'b11000100010011000000; // C44C0 RSHW
      11'h1CB : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h1CC : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h1CD : r_q_a <= 20'b10100101011010000000; // A5680 LDW DL[EA1].
      11'h1CE : r_q_a <= 20'b01100101000000000000; // 65000 FLAG -----,CIN=T[15]
      11'h1CF : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h1D0 : r_q_a <= 20'b11000101010000110001; // C5431 EXTW
      11'h1D1 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h1D2 : r_q_a <= 20'b10110011010101000000; // B3540 STW DH[EA1]; RTS
      11'h1D3 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h1D4 : r_q_a <= 20'b11000000001001011000; // C0258 TSTB.
      11'h1D5 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h1D6 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h1D7 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h1D8 : r_q_a <= 20'b11000000011001011000; // C0658 TSTW.
      11'h1D9 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h1DA : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h1DB : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h1DC : r_q_a <= 20'b11000000011001011000; // C0658 TSTW.
      11'h1DD : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h1DE : r_q_a <= 20'b11000000101001011000; // C0A58 TSTL.
      11'h1DF : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h1E0 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h1E1 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h1E2 : r_q_a <= 20'b11000000001001011000; // C0258 TSTB.
      11'h1E3 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h1E4 : r_q_a <= 20'b01000000000010000000; // 40080 LIT #0080
      11'h1E5 : r_q_a <= 20'b11000011000001011010; // C305A ORB
      11'h1E6 : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h1E7 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h1E8 : r_q_a <= 20'b00101110011000110000; // 2E630 CALL EA1_Calc
      11'h1E9 : r_q_a <= 20'b00000000000111110000; // 001F0 LOOP #16
      11'h1EA : r_q_a <= 20'b00110100100111110000; // 349F0 JUMPN T[0],NoMoveW_r
      11'h1EB : r_q_a <= 20'b10000101010110000100; // 85584 LDW (EA1)+
      11'h1EC : r_q_a <= 20'b01100101000000000000; // 65000 FLAG -----,CIN=T[15]
      11'h1ED : r_q_a <= 20'b10100011010001000111; // A3447 STW RL[CNT]
      11'h1EE : r_q_a <= 20'b11000101010000110001; // C5431 EXTW
      11'h1EF : r_q_a <= 20'b10100011010101000111; // A3547 STW RH[CNT]
      11'h1F0 : r_q_a <= 20'b11000100010011000000; // C44C0 RSHW
      11'h1F1 : r_q_a <= 20'b01100000100000000000; // 60800 FLAG -----,CIN=CLR
      11'h1F2 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h1F3 : r_q_a <= 20'b00101110000111100111; // 2E1E7 CALL Op_MOVEMW_r
      11'h1F4 : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h1F5 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h1F6 : r_q_a <= 20'b00101110011000110000; // 2E630 CALL EA1_Calc
      11'h1F7 : r_q_a <= 20'b00000000000111111101; // 001FD LOOP #16
      11'h1F8 : r_q_a <= 20'b00110100100111111101; // 349FD JUMPN T[0],NoMoveL_r
      11'h1F9 : r_q_a <= 20'b10000101010110000100; // 85584 LDW (EA1)+
      11'h1FA : r_q_a <= 20'b10100011010101000111; // A3547 STW RH[CNT]
      11'h1FB : r_q_a <= 20'b10000101010110000100; // 85584 LDW (EA1)+
      11'h1FC : r_q_a <= 20'b10100011010001000111; // A3447 STW RL[CNT]
      11'h1FD : r_q_a <= 20'b11000100010011000000; // C44C0 RSHW
      11'h1FE : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h1FF : r_q_a <= 20'b00101110000111110101; // 2E1F5 CALL Op_MOVEML_r
      11'h200 : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h201 : r_q_a <= 20'b11010000010001011000; // D0458 NOP; RTS
      11'h202 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h203 : r_q_a <= 20'b00111110000001000001; // 3E041 JUMP Trap_Processing
      11'h204 : r_q_a <= 20'b10000000010110001010; // 8058A FTW (PC)+
      11'h205 : r_q_a <= 20'b00101110011010110010; // 2E6B2 CALL SP_to_EA2
      11'h206 : r_q_a <= 20'b10100101010110000001; // A5581 LDW AH[EA1]
      11'h207 : r_q_a <= 20'b10100101010010000001; // A5481 LDW AL[EA1]
      11'h208 : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h209 : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h20A : r_q_a <= 20'b10000101010010000011; // 85483 LDW EA2H
      11'h20B : r_q_a <= 20'b10100000010101000001; // A0541 WRW AH[EA1]
      11'h20C : r_q_a <= 20'b10000101010010000010; // 85482 LDW EA2L
      11'h20D : r_q_a <= 20'b10100000010001000001; // A0441 WRW AL[EA1]
      11'h20E : r_q_a <= 20'b00101110011010001111; // 2E68F CALL AddOffs
      11'h20F : r_q_a <= 20'b10100011010101000011; // A3543 STW A7H
      11'h210 : r_q_a <= 20'b10110011010001000011; // B3443 STW A7L; RTS
      11'h211 : r_q_a <= 20'b10100101010110000001; // A5581 LDW AH[EA1]
      11'h212 : r_q_a <= 20'b10000011010001000011; // 83443 STW EA2H
      11'h213 : r_q_a <= 20'b10100101010010000001; // A5481 LDW AL[EA1]
      11'h214 : r_q_a <= 20'b10000011010001000010; // 83442 STW EA2L
      11'h215 : r_q_a <= 20'b10000101010110000101; // 85585 LDW (EA2)+
      11'h216 : r_q_a <= 20'b10100011010101000001; // A3541 STW AH[EA1]
      11'h217 : r_q_a <= 20'b10000101010110000101; // 85585 LDW (EA2)+
      11'h218 : r_q_a <= 20'b10100011010001000001; // A3441 STW AL[EA1]
      11'h219 : r_q_a <= 20'b10000101010010000011; // 85483 LDW EA2H
      11'h21A : r_q_a <= 20'b10100011010101000011; // A3543 STW A7H
      11'h21B : r_q_a <= 20'b10000101010010000010; // 85482 LDW EA2L
      11'h21C : r_q_a <= 20'b10110011010001000011; // B3443 STW A7L; RTS
      11'h21D : r_q_a <= 20'b10100101010110000001; // A5581 LDW AH[EA1]
      11'h21E : r_q_a <= 20'b10100101010010000001; // A5481 LDW AL[EA1]
      11'h21F : r_q_a <= 20'b10100011010001001110; // A344E STW USPL
      11'h220 : r_q_a <= 20'b10110011010101001110; // B354E STW USPH; RTS
      11'h221 : r_q_a <= 20'b10100101010110001110; // A558E LDW USPH
      11'h222 : r_q_a <= 20'b10100101010010001110; // A548E LDW USPL
      11'h223 : r_q_a <= 20'b10100011010001000001; // A3441 STW AL[EA1]
      11'h224 : r_q_a <= 20'b10110011010101000001; // B3541 STW AH[EA1]; RTS
      11'h225 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h226 : r_q_a <= 20'b10000011010001001111; // 8344F STW SR
      11'h227 : r_q_a <= 20'b00111011101000100111; // 3BA27 JUMPN I_SR,Op_STOP_Wait
      11'h228 : r_q_a <= 20'b00111110011011001000; // 3E6C8 JUMP Leave_Super
      11'h229 : r_q_a <= 20'b00101110011010110010; // 2E6B2 CALL SP_to_EA2
      11'h22A : r_q_a <= 20'b10000101010110000101; // 85585 LDW (EA2)+
      11'h22B : r_q_a <= 20'b10000011010001001111; // 8344F STW SR
      11'h22C : r_q_a <= 20'b00101110001000101111; // 2E22F CALL Op_RTS_jmp
      11'h22D : r_q_a <= 20'b00111110011011001000; // 3E6C8 JUMP Leave_Super
      11'h22E : r_q_a <= 20'b00101110011010110010; // 2E6B2 CALL SP_to_EA2
      11'h22F : r_q_a <= 20'b10000101010110000101; // 85585 LDW (EA2)+
      11'h230 : r_q_a <= 20'b10000011010001000101; // 83445 STW PCH
      11'h231 : r_q_a <= 20'b10000101010110000101; // 85585 LDW (EA2)+
      11'h232 : r_q_a <= 20'b10000011010001000100; // 83444 STW PCL
      11'h233 : r_q_a <= 20'b00111110011010101110; // 3E6AE JUMP EA2_to_SP
      11'h234 : r_q_a <= 20'b00111000101000000001; // 38A01 JUMPN V_SR,Op_NOP
      11'h235 : r_q_a <= 20'b01000000000000011100; // 4001C LIT #001C
      11'h236 : r_q_a <= 20'b00111110000001000001; // 3E041 JUMP Trap_Processing
      11'h237 : r_q_a <= 20'b00101110011010110010; // 2E6B2 CALL SP_to_EA2
      11'h238 : r_q_a <= 20'b10000101010110000101; // 85585 LDW (EA2)+
      11'h239 : r_q_a <= 20'b10000011000001001111; // 8304F STB SR
      11'h23A : r_q_a <= 20'b00111110001000101111; // 3E22F JUMP Op_RTS_jmp
      11'h23B : r_q_a <= 20'b00101110011000110000; // 2E630 CALL EA1_Calc
      11'h23C : r_q_a <= 20'b00101110011010101001; // 2E6A9 CALL PC_to_Stack
      11'h23D : r_q_a <= 20'b10000101010010000001; // 85481 LDW EA1H
      11'h23E : r_q_a <= 20'b10000011010001000101; // 83445 STW PCH
      11'h23F : r_q_a <= 20'b10000101010010000000; // 85480 LDW EA1L
      11'h240 : r_q_a <= 20'b10010011010001000100; // 93444 STW PCL; RTS
      11'h241 : r_q_a <= 20'b00101110011000110000; // 2E630 CALL EA1_Calc
      11'h242 : r_q_a <= 20'b00111110001000111101; // 3E23D JUMP EA1_to_PC
      11'h243 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h244 : r_q_a <= 20'b10100101011010000100; // A5684 LDW DL[EA2].
      11'h245 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h246 : r_q_a <= 20'b00111001001001001110; // 3924E JUMP N_SR,Trap_Neg
      11'h247 : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h248 : r_q_a <= 20'b00110011001001001010; // 3324A JUMP G_FLG,Trap_Grt
      11'h249 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h24A : r_q_a <= 20'b01100000100100000000; // 60900 FLAG -0---,CIN=CLR
      11'h24B : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h24C : r_q_a <= 20'b01000000000000011000; // 40018 LIT #0018
      11'h24D : r_q_a <= 20'b00111110000001000001; // 3E041 JUMP Trap_Processing
      11'h24E : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h24F : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h250 : r_q_a <= 20'b01000000000000011000; // 40018 LIT #0018
      11'h251 : r_q_a <= 20'b00111110000001000001; // 3E041 JUMP Trap_Processing
      11'h252 : r_q_a <= 20'b00101110011000110000; // 2E630 CALL EA1_Calc
      11'h253 : r_q_a <= 20'b10000101010010000000; // 85480 LDW EA1L
      11'h254 : r_q_a <= 20'b10100011010001000101; // A3445 STW AL[EA2]
      11'h255 : r_q_a <= 20'b10000101010010000001; // 85481 LDW EA1H
      11'h256 : r_q_a <= 20'b10110011010101000101; // B3545 STW AH[EA2]; RTS
      11'h257 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h258 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h259 : r_q_a <= 20'b11000011001000001010; // C320A ADDB.
      11'h25A : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h25B : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h25C : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h25D : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h25E : r_q_a <= 20'b11000011011000001010; // C360A ADDW.
      11'h25F : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h260 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h261 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h262 : r_q_a <= 20'b10100011010001001100; // A344C STW TMP1L
      11'h263 : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h264 : r_q_a <= 20'b10100101010010001100; // A548C LDW TMP1L
      11'h265 : r_q_a <= 20'b11000011011000001010; // C360A ADDW.
      11'h266 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h267 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h268 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h269 : r_q_a <= 20'b11000011101000011010; // C3A1A ADDCL.
      11'h26A : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h26B : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h26C : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h26D : r_q_a <= 20'b10100101010010000001; // A5481 LDW AL[EA1]
      11'h26E : r_q_a <= 20'b11000011011000001010; // C360A ADDW.
      11'h26F : r_q_a <= 20'b10100011010001000001; // A3441 STW AL[EA1]
      11'h270 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h271 : r_q_a <= 20'b10100101010110000001; // A5581 LDW AH[EA1]
      11'h272 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h273 : r_q_a <= 20'b11000011101000011010; // C3A1A ADDCL.
      11'h274 : r_q_a <= 20'b10110011010101000001; // B3541 STW AH[EA1]; RTS
      11'h275 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h276 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h277 : r_q_a <= 20'b11000011001000101011; // C322B SUBB.
      11'h278 : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h279 : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h27A : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h27B : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h27C : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h27D : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h27E : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h27F : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h280 : r_q_a <= 20'b10100011010001001100; // A344C STW TMP1L
      11'h281 : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h282 : r_q_a <= 20'b10100101010010001100; // A548C LDW TMP1L
      11'h283 : r_q_a <= 20'b11000011011000101110; // C362E SUBW.
      11'h284 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h285 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h286 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h287 : r_q_a <= 20'b11000011101000111110; // C3A3E SUBCL.
      11'h288 : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h289 : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h28A : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h28B : r_q_a <= 20'b10100101010010000001; // A5481 LDW AL[EA1]
      11'h28C : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h28D : r_q_a <= 20'b10100011010001000001; // A3441 STW AL[EA1]
      11'h28E : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h28F : r_q_a <= 20'b10100101010110000001; // A5581 LDW AH[EA1]
      11'h290 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h291 : r_q_a <= 20'b11000011101000111011; // C3A3B SUBCL.
      11'h292 : r_q_a <= 20'b10110011010101000001; // B3541 STW AH[EA1]; RTS
      11'h293 : r_q_a <= 20'b00111010001010010110; // 3A296 JUMP B_SR,Op_Scc_Set
      11'h294 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h295 : r_q_a <= 20'b00111110011000111101; // 3E63D JUMP EA1_Write_B
      11'h296 : r_q_a <= 20'b01000000000011111111; // 400FF LIT #00FF
      11'h297 : r_q_a <= 20'b00111110011000111101; // 3E63D JUMP EA1_Write_B
      11'h298 : r_q_a <= 20'b00111010101010011010; // 3AA9A JUMPN B_SR,Op_DBcc_Exec
      11'h299 : r_q_a <= 20'b10010000010110001010; // 9058A FTW (PC)+; RTS
      11'h29A : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h29B : r_q_a <= 20'b11000000010000001001; // C0409 DECW
      11'h29C : r_q_a <= 20'b10100000010001000000; // A0440 WRW DL[EA1]
      11'h29D : r_q_a <= 20'b11000000011001111010; // C067A NOTW.
      11'h29E : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h29F : r_q_a <= 20'b00110001001010011001; // 31299 JUMP Z_FLG,Op_DBcc_Exit
      11'h2A0 : r_q_a <= 20'b10000101010010000101; // 85485 LDW PCH
      11'h2A1 : r_q_a <= 20'b10000101010010000100; // 85484 LDW PCL
      11'h2A2 : r_q_a <= 20'b10000000010110001010; // 8058A FTW (PC)+
      11'h2A3 : r_q_a <= 20'b00111110001010101000; // 3E2A8 JUMP AddWOffs_PC
      11'h2A4 : r_q_a <= 20'b00111010101010110000; // 3AAB0 JUMPN B_SR,FetchDisp
      11'h2A5 : r_q_a <= 20'b10000101010010000101; // 85485 LDW PCH
      11'h2A6 : r_q_a <= 20'b10000101010010000100; // 85484 LDW PCL
      11'h2A7 : r_q_a <= 20'b00101110001010110000; // 2E2B0 CALL FetchDisp
      11'h2A8 : r_q_a <= 20'b00101110011010001111; // 2E68F CALL AddOffs
      11'h2A9 : r_q_a <= 20'b10000011010001000101; // 83445 STW PCH
      11'h2AA : r_q_a <= 20'b10010011010001000100; // 93444 STW PCL; RTS
      11'h2AB : r_q_a <= 20'b10000101010010000101; // 85485 LDW PCH
      11'h2AC : r_q_a <= 20'b10000101010010000100; // 85484 LDW PCL
      11'h2AD : r_q_a <= 20'b00101110001010110000; // 2E2B0 CALL FetchDisp
      11'h2AE : r_q_a <= 20'b00101110011010101001; // 2E6A9 CALL PC_to_Stack
      11'h2AF : r_q_a <= 20'b00111110001010101000; // 3E2A8 JUMP AddWOffs_PC
      11'h2B0 : r_q_a <= 20'b10000101011010001000; // 85688 LDW IMM.
      11'h2B1 : r_q_a <= 20'b00110001101010110100; // 31AB4 JUMPN Z_FLG,ShortBranch
      11'h2B2 : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h2B3 : r_q_a <= 20'b10010000010110001010; // 9058A FTW (PC)+; RTS
      11'h2B4 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h2B5 : r_q_a <= 20'b10000101011010001000; // 85688 LDW IMM.
      11'h2B6 : r_q_a <= 20'b01100101000000000000; // 65000 FLAG -----,CIN=T[15]
      11'h2B7 : r_q_a <= 20'b11000101010000110001; // C5431 EXTW
      11'h2B8 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h2B9 : r_q_a <= 20'b10100011010101000100; // A3544 STW DH[EA2]
      11'h2BA : r_q_a <= 20'b10110011010001000100; // B3444 STW DL[EA2]; RTS
      11'h2BB : r_q_a <= 20'b00101110001010111111; // 2E2BF CALL Op_ORB
      11'h2BC : r_q_a <= 20'b10110011000001000100; // B3044 STB DL[EA2]; RTS
      11'h2BD : r_q_a <= 20'b00101110001010111111; // 2E2BF CALL Op_ORB
      11'h2BE : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h2BF : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h2C0 : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h2C1 : r_q_a <= 20'b11000011001001011010; // C325A ORB.
      11'h2C2 : r_q_a <= 20'b01110000100010011010; // 7089A FLAG -**00,CIN=CLR; RTS
      11'h2C3 : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h2C4 : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h2C5 : r_q_a <= 20'b00101110001011001101; // 2E2CD CALL SBCD_Calc
      11'h2C6 : r_q_a <= 20'b01100000100011010000; // 608D0 FLAG -*#--,CIN=CLR
      11'h2C7 : r_q_a <= 20'b10110011000001000100; // B3044 STB DL[EA2]; RTS
      11'h2C8 : r_q_a <= 20'b00101110011100111101; // 2E73D CALL EA1_RB_An_Dec
      11'h2C9 : r_q_a <= 20'b00101110011001100001; // 2E661 CALL EA2_RB_An_Dec
      11'h2CA : r_q_a <= 20'b00101110001011001101; // 2E2CD CALL SBCD_Calc
      11'h2CB : r_q_a <= 20'b01100000100011010000; // 608D0 FLAG -*#--,CIN=CLR
      11'h2CC : r_q_a <= 20'b10010011000101000101; // 93145 STB (EA2)+; RTS
      11'h2CD : r_q_a <= 20'b11000101010001010010; // C5452 OVER
      11'h2CE : r_q_a <= 20'b01000000000000001111; // 4000F LIT #000F
      11'h2CF : r_q_a <= 20'b11000011010001001010; // C344A ANDW
      11'h2D0 : r_q_a <= 20'b11000101010001010010; // C5452 OVER
      11'h2D1 : r_q_a <= 20'b01000000000000001111; // 4000F LIT #000F
      11'h2D2 : r_q_a <= 20'b11000011010001001010; // C344A ANDW
      11'h2D3 : r_q_a <= 20'b01100010010000000010; // 62402 FLAG 0---0,CIN=X_SR
      11'h2D4 : r_q_a <= 20'b11000011011000111011; // C363B SUBCW.
      11'h2D5 : r_q_a <= 20'b00110010101011011000; // 32AD8 JUMPN N_FLG,SBCD_PosLoNib
      11'h2D6 : r_q_a <= 20'b01000000000000000110; // 40006 LIT #0006
      11'h2D7 : r_q_a <= 20'b11000011010000101110; // C342E SUBW
      11'h2D8 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h2D9 : r_q_a <= 20'b01000000000011110000; // 400F0 LIT #00F0
      11'h2DA : r_q_a <= 20'b11000011010001001010; // C344A ANDW
      11'h2DB : r_q_a <= 20'b11000011010000001010; // C340A ADDW
      11'h2DC : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h2DD : r_q_a <= 20'b01000000000011110000; // 400F0 LIT #00F0
      11'h2DE : r_q_a <= 20'b11000011010001001010; // C344A ANDW
      11'h2DF : r_q_a <= 20'b11000011011000101110; // C362E SUBW.
      11'h2E0 : r_q_a <= 20'b00110010101011100100; // 32AE4 JUMPN N_FLG,SBCD_PosHiNib
      11'h2E1 : r_q_a <= 20'b01000000000001100000; // 40060 LIT #0060
      11'h2E2 : r_q_a <= 20'b11000011010000101110; // C342E SUBW
      11'h2E3 : r_q_a <= 20'b01100000011000000011; // 60603 FLAG 1---1,CIN=KEEP
      11'h2E4 : r_q_a <= 20'b11010000011001011000; // D0658 NOP.; RTS
      11'h2E5 : r_q_a <= 20'b00101110001011101001; // 2E2E9 CALL Op_ORW
      11'h2E6 : r_q_a <= 20'b10110011010001000100; // B3444 STW DL[EA2]; RTS
      11'h2E7 : r_q_a <= 20'b00101110001011101001; // 2E2E9 CALL Op_ORW
      11'h2E8 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h2E9 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h2EA : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h2EB : r_q_a <= 20'b11000011011001011010; // C365A ORW.
      11'h2EC : r_q_a <= 20'b01110000100010011010; // 7089A FLAG -**00,CIN=CLR; RTS
      11'h2ED : r_q_a <= 20'b00101110001011110001; // 2E2F1 CALL Op_ORL
      11'h2EE : r_q_a <= 20'b00111110011010000010; // 3E682 JUMP EA2_WL_Reg
      11'h2EF : r_q_a <= 20'b00101110001011110001; // 2E2F1 CALL Op_ORL
      11'h2F0 : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h2F1 : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h2F2 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h2F3 : r_q_a <= 20'b11000011011001011010; // C365A ORW.
      11'h2F4 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h2F5 : r_q_a <= 20'b10100101010110000100; // A5584 LDW DH[EA2]
      11'h2F6 : r_q_a <= 20'b11000011101001011010; // C3A5A ORL.
      11'h2F7 : r_q_a <= 20'b01110000100010011010; // 7089A FLAG -**00,CIN=CLR; RTS
      11'h2F8 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h2F9 : r_q_a <= 20'b01100000100000000010; // 60802 FLAG ----0,CIN=CLR
      11'h2FA : r_q_a <= 20'b11000000011001011000; // C0658 TSTW.
      11'h2FB : r_q_a <= 20'b00110001000000110110; // 31036 JUMP Z_FLG,Trap_DivZero
      11'h2FC : r_q_a <= 20'b10100101010110000100; // A5584 LDW DH[EA2]
      11'h2FD : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h2FE : r_q_a <= 20'b00101110001100000011; // 2E303 CALL Op_DIVx
      11'h2FF : r_q_a <= 20'b00111000001100010011; // 38313 JUMP V_SR,Op_Div_Overflow2
      11'h300 : r_q_a <= 20'b01100000100010010010; // 60892 FLAG -**-0,CIN=CLR
      11'h301 : r_q_a <= 20'b10100011010001000100; // A3444 STW DL[EA2]
      11'h302 : r_q_a <= 20'b10110011010101000100; // B3544 STW DH[EA2]; RTS
      11'h303 : r_q_a <= 20'b01100000100000000010; // 60802 FLAG ----0,CIN=CLR
      11'h304 : r_q_a <= 20'b10000011010001001010; // 8344A STW ACCL
      11'h305 : r_q_a <= 20'b10000011010001001011; // 8344B STW ACCH
      11'h306 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h307 : r_q_a <= 20'b10000000010001001001; // 80449 WRW LSHR
      11'h308 : r_q_a <= 20'b11000100101011100000; // C4AE0 DIV.
      11'h309 : r_q_a <= 20'b00000000001100001010; // 0030A LOOP #16
      11'h30A : r_q_a <= 20'b11000100101011100000; // C4AE0 DIV.
      11'h30B : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h30C : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h30D : r_q_a <= 20'b01100000100000000100; // 60804 FLAG ---*-,CIN=CLR
      11'h30E : r_q_a <= 20'b00111000001100010011; // 38313 JUMP V_SR,Op_Div_Overflow2
      11'h30F : r_q_a <= 20'b10000101010010001010; // 8548A LDW ACCL
      11'h310 : r_q_a <= 20'b10010101011010001001; // 95689 LDW LSHR.; RTS
      11'h311 : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h312 : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h313 : r_q_a <= 20'b01110000100000001100; // 7080C FLAG ---1-,CIN=CLR; RTS
      11'h314 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h315 : r_q_a <= 20'b01100000100000000010; // 60802 FLAG ----0,CIN=CLR
      11'h316 : r_q_a <= 20'b11000000011001011000; // C0658 TSTW.
      11'h317 : r_q_a <= 20'b00110001000000110110; // 31036 JUMP Z_FLG,Trap_DivZero
      11'h318 : r_q_a <= 20'b00110010101100101000; // 32B28 JUMPN N_FLG,Op_DIVS_Src_Pos
      11'h319 : r_q_a <= 20'b11000000010000101100; // C042C NEGW
      11'h31A : r_q_a <= 20'b10100101011110000100; // A5784 LDW DH[EA2].
      11'h31B : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h31C : r_q_a <= 20'b00110010101100110000; // 32B30 JUMPN N_FLG,Op_DIVS_Neg
      11'h31D : r_q_a <= 20'b11000000011000101100; // C062C NEGW.
      11'h31E : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h31F : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h320 : r_q_a <= 20'b11000000101000111100; // C0A3C NEGCL.
      11'h321 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h322 : r_q_a <= 20'b00101110001100000011; // 2E303 CALL Op_DIVx
      11'h323 : r_q_a <= 20'b00111000001100010011; // 38313 JUMP V_SR,Op_Div_Overflow2
      11'h324 : r_q_a <= 20'b00110010001100010001; // 32311 JUMP N_FLG,Op_Div_Overflow
      11'h325 : r_q_a <= 20'b01100000100010010010; // 60892 FLAG -**-0,CIN=CLR
      11'h326 : r_q_a <= 20'b10100011010001000100; // A3444 STW DL[EA2]
      11'h327 : r_q_a <= 20'b10110011010101000100; // B3544 STW DH[EA2]; RTS
      11'h328 : r_q_a <= 20'b10100101011110000100; // A5784 LDW DH[EA2].
      11'h329 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h32A : r_q_a <= 20'b00110010101100100010; // 32B22 JUMPN N_FLG,Op_DIVS_Pos
      11'h32B : r_q_a <= 20'b11000000011000101100; // C062C NEGW.
      11'h32C : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h32D : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h32E : r_q_a <= 20'b11000000101000111100; // C0A3C NEGCL.
      11'h32F : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h330 : r_q_a <= 20'b00101110001100000011; // 2E303 CALL Op_DIVx
      11'h331 : r_q_a <= 20'b00111000001100010011; // 38313 JUMP V_SR,Op_Div_Overflow2
      11'h332 : r_q_a <= 20'b00110010001100010001; // 32311 JUMP N_FLG,Op_Div_Overflow
      11'h333 : r_q_a <= 20'b11000000011000101100; // C062C NEGW.
      11'h334 : r_q_a <= 20'b01100000100010010010; // 60892 FLAG -**-0,CIN=CLR
      11'h335 : r_q_a <= 20'b10100011010001000100; // A3444 STW DL[EA2]
      11'h336 : r_q_a <= 20'b10110011010101000100; // B3544 STW DH[EA2]; RTS
      11'h337 : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h338 : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h339 : r_q_a <= 20'b11000011001000101011; // C322B SUBB.
      11'h33A : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h33B : r_q_a <= 20'b10110011000001000100; // B3044 STB DL[EA2]; RTS
      11'h33C : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h33D : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h33E : r_q_a <= 20'b11000011001000101011; // C322B SUBB.
      11'h33F : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h340 : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h341 : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h342 : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h343 : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h344 : r_q_a <= 20'b11000011001000111011; // C323B SUBCB.
      11'h345 : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h346 : r_q_a <= 20'b10110011000001000100; // B3044 STB DL[EA2]; RTS
      11'h347 : r_q_a <= 20'b00101110011100111101; // 2E73D CALL EA1_RB_An_Dec
      11'h348 : r_q_a <= 20'b00101110011001100001; // 2E661 CALL EA2_RB_An_Dec
      11'h349 : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h34A : r_q_a <= 20'b11000011001000111011; // C323B SUBCB.
      11'h34B : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h34C : r_q_a <= 20'b10010011000101000101; // 93145 STB (EA2)+; RTS
      11'h34D : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h34E : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h34F : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h350 : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h351 : r_q_a <= 20'b10110011010001000100; // B3444 STW DL[EA2]; RTS
      11'h352 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h353 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h354 : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h355 : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h356 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h357 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h358 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h359 : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h35A : r_q_a <= 20'b11000011011000111011; // C363B SUBCW.
      11'h35B : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h35C : r_q_a <= 20'b10110011010001000100; // B3444 STW DL[EA2]; RTS
      11'h35D : r_q_a <= 20'b00101110011101001101; // 2E74D CALL EA1_RW_An_Dec
      11'h35E : r_q_a <= 20'b00101110011001100111; // 2E667 CALL EA2_RW_An_Dec
      11'h35F : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h360 : r_q_a <= 20'b11000011011000111011; // C363B SUBCW.
      11'h361 : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h362 : r_q_a <= 20'b10010011010101000001; // 93541 STW (EA2); RTS
      11'h363 : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h364 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h365 : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h366 : r_q_a <= 20'b10100011010001000100; // A3444 STW DL[EA2]
      11'h367 : r_q_a <= 20'b10100101010110000100; // A5584 LDW DH[EA2]
      11'h368 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h369 : r_q_a <= 20'b11000011101000111011; // C3A3B SUBCL.
      11'h36A : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h36B : r_q_a <= 20'b10110011010101000100; // B3544 STW DH[EA2]; RTS
      11'h36C : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h36D : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h36E : r_q_a <= 20'b11000011011000101110; // C362E SUBW.
      11'h36F : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h370 : r_q_a <= 20'b10100101010110000100; // A5584 LDW DH[EA2]
      11'h371 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h372 : r_q_a <= 20'b11000011101000111110; // C3A3E SUBCL.
      11'h373 : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h374 : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h375 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h376 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h377 : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h378 : r_q_a <= 20'b11000011011000111011; // C363B SUBCW.
      11'h379 : r_q_a <= 20'b10100011010001000100; // A3444 STW DL[EA2]
      11'h37A : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h37B : r_q_a <= 20'b10100101010110000100; // A5584 LDW DH[EA2]
      11'h37C : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h37D : r_q_a <= 20'b11000011101000111011; // C3A3B SUBCL.
      11'h37E : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h37F : r_q_a <= 20'b10110011010101000100; // B3544 STW DH[EA2]; RTS
      11'h380 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h381 : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h382 : r_q_a <= 20'b10000101010110001000; // 85588 LDW -(EA1)
      11'h383 : r_q_a <= 20'b10000101010110001001; // 85589 LDW -(EA2)
      11'h384 : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h385 : r_q_a <= 20'b11000011011000111011; // C363B SUBCW.
      11'h386 : r_q_a <= 20'b10000101010110001000; // 85588 LDW -(EA1)
      11'h387 : r_q_a <= 20'b10000101010110001001; // 85589 LDW -(EA2)
      11'h388 : r_q_a <= 20'b00101110011011011110; // 2E6DE CALL Set_An_EA1
      11'h389 : r_q_a <= 20'b00101110011100001010; // 2E70A CALL Set_An_EA2
      11'h38A : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h38B : r_q_a <= 20'b11000011101000111011; // C3A3B SUBCL.
      11'h38C : r_q_a <= 20'b10000011010101000101; // 83545 STW (EA2)+
      11'h38D : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h38E : r_q_a <= 20'b10010011010101000001; // 93541 STW (EA2); RTS
      11'h38F : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h390 : r_q_a <= 20'b01100101000000000000; // 65000 FLAG -----,CIN=T[15]
      11'h391 : r_q_a <= 20'b11000101010000110001; // C5431 EXTW
      11'h392 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h393 : r_q_a <= 20'b10100101010010000101; // A5485 LDW AL[EA2]
      11'h394 : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h395 : r_q_a <= 20'b10100011010001000101; // A3445 STW AL[EA2]
      11'h396 : r_q_a <= 20'b10100101010110000101; // A5585 LDW AH[EA2]
      11'h397 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h398 : r_q_a <= 20'b11000011100000111011; // C383B SUBCL
      11'h399 : r_q_a <= 20'b10110011010101000101; // B3545 STW AH[EA2]; RTS
      11'h39A : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h39B : r_q_a <= 20'b00111110001110010011; // 3E393 JUMP Op_SUBA_jmp
      11'h39C : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h39D : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h39E : r_q_a <= 20'b11000011001000101011; // C322B SUBB.
      11'h39F : r_q_a <= 20'b01100000100010010101; // 60895 FLAG -****,CIN=CLR
      11'h3A0 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h3A1 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h3A2 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h3A3 : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h3A4 : r_q_a <= 20'b01100000100010010101; // 60895 FLAG -****,CIN=CLR
      11'h3A5 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h3A6 : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h3A7 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h3A8 : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h3A9 : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h3AA : r_q_a <= 20'b10100101010110000100; // A5584 LDW DH[EA2]
      11'h3AB : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h3AC : r_q_a <= 20'b11000011101000111011; // C3A3B SUBCL.
      11'h3AD : r_q_a <= 20'b01100000100010010101; // 60895 FLAG -****,CIN=CLR
      11'h3AE : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h3AF : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h3B0 : r_q_a <= 20'b01100101000000000000; // 65000 FLAG -----,CIN=T[15]
      11'h3B1 : r_q_a <= 20'b11000101010000110001; // C5431 EXTW
      11'h3B2 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h3B3 : r_q_a <= 20'b10100101010010000101; // A5485 LDW AL[EA2]
      11'h3B4 : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h3B5 : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h3B6 : r_q_a <= 20'b10100101010110000101; // A5585 LDW AH[EA2]
      11'h3B7 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h3B8 : r_q_a <= 20'b11000011101000111011; // C3A3B SUBCL.
      11'h3B9 : r_q_a <= 20'b01100000100010010101; // 60895 FLAG -****,CIN=CLR
      11'h3BA : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h3BB : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h3BC : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h3BD : r_q_a <= 20'b11000011001001101010; // C326A XORB.
      11'h3BE : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h3BF : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h3C0 : r_q_a <= 20'b00101110010111110011; // 2E5F3 CALL EA1_RB_An_Inc
      11'h3C1 : r_q_a <= 20'b00101110011001011110; // 2E65E CALL EA2_RB_An_Inc
      11'h3C2 : r_q_a <= 20'b11000011001000101011; // C322B SUBB.
      11'h3C3 : r_q_a <= 20'b01100000100010010101; // 60895 FLAG -****,CIN=CLR
      11'h3C4 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h3C5 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h3C6 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h3C7 : r_q_a <= 20'b11000011011001101010; // C366A XORW.
      11'h3C8 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h3C9 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h3CA : r_q_a <= 20'b00101110011000000100; // 2E604 CALL EA1_RW_An_Inc
      11'h3CB : r_q_a <= 20'b00101110011001100100; // 2E664 CALL EA2_RW_An_Inc
      11'h3CC : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h3CD : r_q_a <= 20'b01100000100010010101; // 60895 FLAG -****,CIN=CLR
      11'h3CE : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h3CF : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h3D0 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h3D1 : r_q_a <= 20'b11000011011001101010; // C366A XORW.
      11'h3D2 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h3D3 : r_q_a <= 20'b10100101010110000100; // A5584 LDW DH[EA2]
      11'h3D4 : r_q_a <= 20'b11000011101001101010; // C3A6A XORL.
      11'h3D5 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h3D6 : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h3D7 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h3D8 : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h3D9 : r_q_a <= 20'b10000101010110000100; // 85584 LDW (EA1)+
      11'h3DA : r_q_a <= 20'b10000101010110000101; // 85585 LDW (EA2)+
      11'h3DB : r_q_a <= 20'b10000101010110000100; // 85584 LDW (EA1)+
      11'h3DC : r_q_a <= 20'b10000101010110000101; // 85585 LDW (EA2)+
      11'h3DD : r_q_a <= 20'b00101110011011011110; // 2E6DE CALL Set_An_EA1
      11'h3DE : r_q_a <= 20'b00101110011100001010; // 2E70A CALL Set_An_EA2
      11'h3DF : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h3E0 : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h3E1 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h3E2 : r_q_a <= 20'b11000011101000111011; // C3A3B SUBCL.
      11'h3E3 : r_q_a <= 20'b01100000100010010101; // 60895 FLAG -****,CIN=CLR
      11'h3E4 : r_q_a <= 20'b11010011010001010010; // D3452 DROP; RTS
      11'h3E5 : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h3E6 : r_q_a <= 20'b00111110001110110011; // 3E3B3 JUMP Op_CMPA
      11'h3E7 : r_q_a <= 20'b00101110001111101011; // 2E3EB CALL Op_ANDB
      11'h3E8 : r_q_a <= 20'b10110011000001000100; // B3044 STB DL[EA2]; RTS
      11'h3E9 : r_q_a <= 20'b00101110001111101011; // 2E3EB CALL Op_ANDB
      11'h3EA : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h3EB : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h3EC : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h3ED : r_q_a <= 20'b11000011001001001010; // C324A ANDB.
      11'h3EE : r_q_a <= 20'b01110000100010011010; // 7089A FLAG -**00,CIN=CLR; RTS
      11'h3EF : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h3F0 : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h3F1 : r_q_a <= 20'b00101110001111111001; // 2E3F9 CALL ABCD_Calc
      11'h3F2 : r_q_a <= 20'b01100000100011010000; // 608D0 FLAG -*#--,CIN=CLR
      11'h3F3 : r_q_a <= 20'b10110011000001000100; // B3044 STB DL[EA2]; RTS
      11'h3F4 : r_q_a <= 20'b00101110011100111101; // 2E73D CALL EA1_RB_An_Dec
      11'h3F5 : r_q_a <= 20'b00101110011001100001; // 2E661 CALL EA2_RB_An_Dec
      11'h3F6 : r_q_a <= 20'b00101110001111111001; // 2E3F9 CALL ABCD_Calc
      11'h3F7 : r_q_a <= 20'b01100000100011010000; // 608D0 FLAG -*#--,CIN=CLR
      11'h3F8 : r_q_a <= 20'b10010011000101000101; // 93145 STB (EA2)+; RTS
      11'h3F9 : r_q_a <= 20'b11000101010001010010; // C5452 OVER
      11'h3FA : r_q_a <= 20'b01000000000000001111; // 4000F LIT #000F
      11'h3FB : r_q_a <= 20'b11000011010001001010; // C344A ANDW
      11'h3FC : r_q_a <= 20'b11000101010001010010; // C5452 OVER
      11'h3FD : r_q_a <= 20'b01000000000000001111; // 4000F LIT #000F
      11'h3FE : r_q_a <= 20'b11000011011001001010; // C364A ANDW.
      11'h3FF : r_q_a <= 20'b01100010010000000010; // 62402 FLAG 0---0,CIN=X_SR
      11'h400 : r_q_a <= 20'b11000011010000011010; // C341A ADDCW
      11'h401 : r_q_a <= 20'b01000000000000001010; // 4000A LIT #000A
      11'h402 : r_q_a <= 20'b11000101010001010010; // C5452 OVER
      11'h403 : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h404 : r_q_a <= 20'b00110010010000001000; // 32408 JUMP N_FLG,ABCD_Less10
      11'h405 : r_q_a <= 20'b01000000000000010000; // 40010 LIT #0010
      11'h406 : r_q_a <= 20'b11000011010000001010; // C340A ADDW
      11'h407 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h408 : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h409 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h40A : r_q_a <= 20'b01000000000011110000; // 400F0 LIT #00F0
      11'h40B : r_q_a <= 20'b11000011010001001010; // C344A ANDW
      11'h40C : r_q_a <= 20'b11000011010000001010; // C340A ADDW
      11'h40D : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h40E : r_q_a <= 20'b01000000000011110000; // 400F0 LIT #00F0
      11'h40F : r_q_a <= 20'b11000011010001001010; // C344A ANDW
      11'h410 : r_q_a <= 20'b11000011010000001010; // C340A ADDW
      11'h411 : r_q_a <= 20'b01000000000010100000; // 400A0 LIT #00A0
      11'h412 : r_q_a <= 20'b11000101010001010010; // C5452 OVER
      11'h413 : r_q_a <= 20'b11000011011000101011; // C362B SUBW.
      11'h414 : r_q_a <= 20'b00110010010000010111; // 32417 JUMP N_FLG,ABCD_Less100
      11'h415 : r_q_a <= 20'b01100000011000000011; // 60603 FLAG 1---1,CIN=KEEP
      11'h416 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h417 : r_q_a <= 20'b11010011011001010010; // D3652 DROP.; RTS
      11'h418 : r_q_a <= 20'b00101110010000011100; // 2E41C CALL Op_ANDW
      11'h419 : r_q_a <= 20'b10110011010001000100; // B3444 STW DL[EA2]; RTS
      11'h41A : r_q_a <= 20'b00101110010000011100; // 2E41C CALL Op_ANDW
      11'h41B : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h41C : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h41D : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h41E : r_q_a <= 20'b11000011011001001010; // C364A ANDW.
      11'h41F : r_q_a <= 20'b01110000100010011010; // 7089A FLAG -**00,CIN=CLR; RTS
      11'h420 : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h421 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h422 : r_q_a <= 20'b10100101010110000100; // A5584 LDW DH[EA2]
      11'h423 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h424 : r_q_a <= 20'b10100011010001000000; // A3440 STW DL[EA1]
      11'h425 : r_q_a <= 20'b10100011010101000000; // A3540 STW DH[EA1]
      11'h426 : r_q_a <= 20'b10100011010001000100; // A3444 STW DL[EA2]
      11'h427 : r_q_a <= 20'b10110011010101000100; // B3544 STW DH[EA2]; RTS
      11'h428 : r_q_a <= 20'b10100101010110000001; // A5581 LDW AH[EA1]
      11'h429 : r_q_a <= 20'b10100101010010000001; // A5481 LDW AL[EA1]
      11'h42A : r_q_a <= 20'b10100101010110000101; // A5585 LDW AH[EA2]
      11'h42B : r_q_a <= 20'b10100101010010000101; // A5485 LDW AL[EA2]
      11'h42C : r_q_a <= 20'b10100011010001000001; // A3441 STW AL[EA1]
      11'h42D : r_q_a <= 20'b10100011010101000001; // A3541 STW AH[EA1]
      11'h42E : r_q_a <= 20'b10100011010001000101; // A3445 STW AL[EA2]
      11'h42F : r_q_a <= 20'b10110011010101000101; // B3545 STW AH[EA2]; RTS
      11'h430 : r_q_a <= 20'b00101110010000110100; // 2E434 CALL Op_ANDL
      11'h431 : r_q_a <= 20'b00111110011010000010; // 3E682 JUMP EA2_WL_Reg
      11'h432 : r_q_a <= 20'b00101110010000110100; // 2E434 CALL Op_ANDL
      11'h433 : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h434 : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h435 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h436 : r_q_a <= 20'b11000011011001001010; // C364A ANDW.
      11'h437 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h438 : r_q_a <= 20'b10100101010110000100; // A5584 LDW DH[EA2]
      11'h439 : r_q_a <= 20'b11000011101001001010; // C3A4A ANDL.
      11'h43A : r_q_a <= 20'b01110000100010011010; // 7089A FLAG -**00,CIN=CLR; RTS
      11'h43B : r_q_a <= 20'b10100101010110000001; // A5581 LDW AH[EA1]
      11'h43C : r_q_a <= 20'b10100101010010000001; // A5481 LDW AL[EA1]
      11'h43D : r_q_a <= 20'b10100101010110000100; // A5584 LDW DH[EA2]
      11'h43E : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h43F : r_q_a <= 20'b10100011010001000001; // A3441 STW AL[EA1]
      11'h440 : r_q_a <= 20'b10100011010101000001; // A3541 STW AH[EA1]
      11'h441 : r_q_a <= 20'b10100011010001000100; // A3444 STW DL[EA2]
      11'h442 : r_q_a <= 20'b10110011010101000100; // B3544 STW DH[EA2]; RTS
      11'h443 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h444 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h445 : r_q_a <= 20'b00101110010001001011; // 2E44B CALL Op_MULx
      11'h446 : r_q_a <= 20'b11000000011001011000; // C0658 TSTW.
      11'h447 : r_q_a <= 20'b10100011010001000100; // A3444 STW DL[EA2]
      11'h448 : r_q_a <= 20'b11000000101001011000; // C0A58 TSTL.
      11'h449 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h44A : r_q_a <= 20'b10110011010101000100; // B3544 STW DH[EA2]; RTS
      11'h44B : r_q_a <= 20'b10000011010001001001; // 83449 STW LSHR
      11'h44C : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h44D : r_q_a <= 20'b10000000010001001010; // 8044A WRW ACCL
      11'h44E : r_q_a <= 20'b10000000010001001011; // 8044B WRW ACCH
      11'h44F : r_q_a <= 20'b01100000100000000000; // 60800 FLAG -----,CIN=CLR
      11'h450 : r_q_a <= 20'b11000100100011000000; // C48C0 RSHL
      11'h451 : r_q_a <= 20'b00000000010001010010; // 00452 LOOP #16
      11'h452 : r_q_a <= 20'b11000100100011110000; // C48F0 MUL
      11'h453 : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h454 : r_q_a <= 20'b11000011010001010010; // C3452 DROP
      11'h455 : r_q_a <= 20'b10000101010010001011; // 8548B LDW ACCH
      11'h456 : r_q_a <= 20'b10010101010010001010; // 9548A LDW ACCL; RTS
      11'h457 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h458 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h459 : r_q_a <= 20'b11000000011001011000; // C0658 TSTW.
      11'h45A : r_q_a <= 20'b00110010110001100000; // 32C60 JUMPN N_FLG,Op_MULS_Src_Pos
      11'h45B : r_q_a <= 20'b11000000010000101100; // C042C NEGW
      11'h45C : r_q_a <= 20'b11000100011001010010; // C4652 SWAP.
      11'h45D : r_q_a <= 20'b00110010110001100011; // 32C63 JUMPN N_FLG,Op_MULS_Neg
      11'h45E : r_q_a <= 20'b11000000010000101100; // C042C NEGW
      11'h45F : r_q_a <= 20'b00111110010001000101; // 3E445 JUMP Op_MULS_Pos
      11'h460 : r_q_a <= 20'b11000100011001010010; // C4652 SWAP.
      11'h461 : r_q_a <= 20'b00110010110001000101; // 32C45 JUMPN N_FLG,Op_MULS_Pos
      11'h462 : r_q_a <= 20'b11000000010000101100; // C042C NEGW
      11'h463 : r_q_a <= 20'b00101110010001001011; // 2E44B CALL Op_MULx
      11'h464 : r_q_a <= 20'b11000000011000101100; // C062C NEGW.
      11'h465 : r_q_a <= 20'b10100011010001000100; // A3444 STW DL[EA2]
      11'h466 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h467 : r_q_a <= 20'b11000000101000111100; // C0A3C NEGCL.
      11'h468 : r_q_a <= 20'b01100000100010011010; // 6089A FLAG -**00,CIN=CLR
      11'h469 : r_q_a <= 20'b10110011010101000100; // B3544 STW DH[EA2]; RTS
      11'h46A : r_q_a <= 20'b00101110010001101110; // 2E46E CALL Op_ADDB
      11'h46B : r_q_a <= 20'b10110011000001000100; // B3044 STB DL[EA2]; RTS
      11'h46C : r_q_a <= 20'b00101110010001101110; // 2E46E CALL Op_ADDB
      11'h46D : r_q_a <= 20'b00111110011000110010; // 3E632 JUMP EA1_Update_B
      11'h46E : r_q_a <= 20'b00101110010111101111; // 2E5EF CALL EA1_Read_B
      11'h46F : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h470 : r_q_a <= 20'b11000011001000001010; // C320A ADDB.
      11'h471 : r_q_a <= 20'b01110000101010010101; // 70A95 FLAG *****,CIN=CLR; RTS
      11'h472 : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h473 : r_q_a <= 20'b10100101000010000100; // A5084 LDB DL[EA2]
      11'h474 : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h475 : r_q_a <= 20'b11000011001000011010; // C321A ADDCB.
      11'h476 : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h477 : r_q_a <= 20'b10110011000001000100; // B3044 STB DL[EA2]; RTS
      11'h478 : r_q_a <= 20'b00101110011100111101; // 2E73D CALL EA1_RB_An_Dec
      11'h479 : r_q_a <= 20'b00101110011001100001; // 2E661 CALL EA2_RB_An_Dec
      11'h47A : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h47B : r_q_a <= 20'b11000011001000011010; // C321A ADDCB.
      11'h47C : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h47D : r_q_a <= 20'b10010011000101000101; // 93145 STB (EA2)+; RTS
      11'h47E : r_q_a <= 20'b00101110010010000010; // 2E482 CALL Op_ADDW
      11'h47F : r_q_a <= 20'b10110011010001000100; // B3444 STW DL[EA2]; RTS
      11'h480 : r_q_a <= 20'b00101110010010000010; // 2E482 CALL Op_ADDW
      11'h481 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h482 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h483 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h484 : r_q_a <= 20'b11000011011000001010; // C360A ADDW.
      11'h485 : r_q_a <= 20'b01110000101010010101; // 70A95 FLAG *****,CIN=CLR; RTS
      11'h486 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h487 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h488 : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h489 : r_q_a <= 20'b11000011011000011010; // C361A ADDCW.
      11'h48A : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h48B : r_q_a <= 20'b10110011010001000100; // B3444 STW DL[EA2]; RTS
      11'h48C : r_q_a <= 20'b00101110011101001101; // 2E74D CALL EA1_RW_An_Dec
      11'h48D : r_q_a <= 20'b00101110011001100111; // 2E667 CALL EA2_RW_An_Dec
      11'h48E : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h48F : r_q_a <= 20'b11000011011000011010; // C361A ADDCW.
      11'h490 : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h491 : r_q_a <= 20'b10010011010101000001; // 93541 STW (EA2); RTS
      11'h492 : r_q_a <= 20'b00101110010010010110; // 2E496 CALL Op_ADDL
      11'h493 : r_q_a <= 20'b00111110011010000010; // 3E682 JUMP EA2_WL_Reg
      11'h494 : r_q_a <= 20'b00101110010010010110; // 2E496 CALL Op_ADDL
      11'h495 : r_q_a <= 20'b00111110011000111010; // 3E63A JUMP EA1_Update_L
      11'h496 : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h497 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h498 : r_q_a <= 20'b11000011011000001010; // C360A ADDW.
      11'h499 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h49A : r_q_a <= 20'b10100101010110000100; // A5584 LDW DH[EA2]
      11'h49B : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h49C : r_q_a <= 20'b11000011101000011010; // C3A1A ADDCL.
      11'h49D : r_q_a <= 20'b01110000101010010101; // 70A95 FLAG *****,CIN=CLR; RTS
      11'h49E : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h49F : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h4A0 : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h4A1 : r_q_a <= 20'b11000011011000011010; // C361A ADDCW.
      11'h4A2 : r_q_a <= 20'b10100011010001000100; // A3444 STW DL[EA2]
      11'h4A3 : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h4A4 : r_q_a <= 20'b10100101010110000100; // A5584 LDW DH[EA2]
      11'h4A5 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h4A6 : r_q_a <= 20'b11000011101000011010; // C3A1A ADDCL.
      11'h4A7 : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h4A8 : r_q_a <= 20'b10110011010101000100; // B3544 STW DH[EA2]; RTS
      11'h4A9 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h4AA : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h4AB : r_q_a <= 20'b10000101010110001000; // 85588 LDW -(EA1)
      11'h4AC : r_q_a <= 20'b10000101010110001001; // 85589 LDW -(EA2)
      11'h4AD : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h4AE : r_q_a <= 20'b11000011011000011010; // C361A ADDCW.
      11'h4AF : r_q_a <= 20'b10000101010110001000; // 85588 LDW -(EA1)
      11'h4B0 : r_q_a <= 20'b10000101010110001001; // 85589 LDW -(EA2)
      11'h4B1 : r_q_a <= 20'b00101110011011011110; // 2E6DE CALL Set_An_EA1
      11'h4B2 : r_q_a <= 20'b00101110011100001010; // 2E70A CALL Set_An_EA2
      11'h4B3 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h4B4 : r_q_a <= 20'b11000011101000011010; // C3A1A ADDCL.
      11'h4B5 : r_q_a <= 20'b10000011010101000101; // 83545 STW (EA2)+
      11'h4B6 : r_q_a <= 20'b01100000101011010101; // 60AD5 FLAG **#**,CIN=CLR
      11'h4B7 : r_q_a <= 20'b10010011010101000001; // 93541 STW (EA2); RTS
      11'h4B8 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h4B9 : r_q_a <= 20'b01100101000000000000; // 65000 FLAG -----,CIN=T[15]
      11'h4BA : r_q_a <= 20'b11000101010000110001; // C5431 EXTW
      11'h4BB : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h4BC : r_q_a <= 20'b10100101010010000101; // A5485 LDW AL[EA2]
      11'h4BD : r_q_a <= 20'b11000011011000001010; // C360A ADDW.
      11'h4BE : r_q_a <= 20'b10100011010001000101; // A3445 STW AL[EA2]
      11'h4BF : r_q_a <= 20'b10100101010110000101; // A5585 LDW AH[EA2]
      11'h4C0 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h4C1 : r_q_a <= 20'b11000011100000011010; // C381A ADDCL
      11'h4C2 : r_q_a <= 20'b10110011010101000101; // B3545 STW AH[EA2]; RTS
      11'h4C3 : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h4C4 : r_q_a <= 20'b00111110010010111100; // 3E4BC JUMP Op_ADDA_jmp
      11'h4C5 : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h4C6 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h4C7 : r_q_a <= 20'b00111110010011001010; // 3E4CA JUMP ASRB_jmp
      11'h4C8 : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h4C9 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h4CA : r_q_a <= 20'b01100110100000001010; // 6680A FLAG ---00,CIN=N[7]
      11'h4CB : r_q_a <= 20'b00000000110011001101; // 00CCD LOOP T
      11'h4CC : r_q_a <= 20'b11000100001011000000; // C42C0 RSHB.
      11'h4CD : r_q_a <= 20'b01100100101000001001; // 64A09 FLAG *--0*,CIN=T[7]
      11'h4CE : r_q_a <= 20'b00111110000110011011; // 3E19B JUMP Write_DnB
      11'h4CF : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h4D0 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h4D1 : r_q_a <= 20'b00111110010011010100; // 3E4D4 JUMP LSRB_jmp
      11'h4D2 : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h4D3 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h4D4 : r_q_a <= 20'b01100000100000001010; // 6080A FLAG ---00,CIN=CLR
      11'h4D5 : r_q_a <= 20'b00000000110011010111; // 00CD7 LOOP T
      11'h4D6 : r_q_a <= 20'b11000100001011000000; // C42C0 RSHB.
      11'h4D7 : r_q_a <= 20'b01100000101000001001; // 60A09 FLAG *--0*,CIN=CLR
      11'h4D8 : r_q_a <= 20'b00111110000110011011; // 3E19B JUMP Write_DnB
      11'h4D9 : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h4DA : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h4DB : r_q_a <= 20'b00111110010011011110; // 3E4DE JUMP ROXRB_jmp
      11'h4DC : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h4DD : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h4DE : r_q_a <= 20'b01100010000000001000; // 62008 FLAG ---0-,CIN=X_SR
      11'h4DF : r_q_a <= 20'b00000000110011100001; // 00CE1 LOOP T
      11'h4E0 : r_q_a <= 20'b11000100001011000000; // C42C0 RSHB.
      11'h4E1 : r_q_a <= 20'b01100001101000001001; // 61A09 FLAG *--0*,CIN=C_FLG
      11'h4E2 : r_q_a <= 20'b00111110000110011011; // 3E19B JUMP Write_DnB
      11'h4E3 : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h4E4 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h4E5 : r_q_a <= 20'b00111110010011101000; // 3E4E8 JUMP RORB_jmp
      11'h4E6 : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h4E7 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h4E8 : r_q_a <= 20'b01100110000000001010; // 6600A FLAG ---00,CIN=N[0]
      11'h4E9 : r_q_a <= 20'b00000000110011101011; // 00CEB LOOP T
      11'h4EA : r_q_a <= 20'b11000100001011000000; // C42C0 RSHB.
      11'h4EB : r_q_a <= 20'b01100100000000001001; // 64009 FLAG ---0*,CIN=T[0]
      11'h4EC : r_q_a <= 20'b00111110000110011011; // 3E19B JUMP Write_DnB
      11'h4ED : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h4EE : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h4EF : r_q_a <= 20'b00111110010011110010; // 3E4F2 JUMP ASLB_jmp
      11'h4F0 : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h4F1 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h4F2 : r_q_a <= 20'b01100000100000001010; // 6080A FLAG ---00,CIN=CLR
      11'h4F3 : r_q_a <= 20'b00000000110011110101; // 00CF5 LOOP T
      11'h4F4 : r_q_a <= 20'b11000100001010000000; // C4280 LSHB.
      11'h4F5 : r_q_a <= 20'b01100000101000000101; // 60A05 FLAG *--**,CIN=CLR
      11'h4F6 : r_q_a <= 20'b00111110000110011011; // 3E19B JUMP Write_DnB
      11'h4F7 : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h4F8 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h4F9 : r_q_a <= 20'b00111110010011111100; // 3E4FC JUMP LSLB_jmp
      11'h4FA : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h4FB : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h4FC : r_q_a <= 20'b01100000100000001010; // 6080A FLAG ---00,CIN=CLR
      11'h4FD : r_q_a <= 20'b00000000110011111111; // 00CFF LOOP T
      11'h4FE : r_q_a <= 20'b11000100001010000000; // C4280 LSHB.
      11'h4FF : r_q_a <= 20'b01100000101000001001; // 60A09 FLAG *--0*,CIN=CLR
      11'h500 : r_q_a <= 20'b00111110000110011011; // 3E19B JUMP Write_DnB
      11'h501 : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h502 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h503 : r_q_a <= 20'b00111110010100000110; // 3E506 JUMP ROXLB_jmp
      11'h504 : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h505 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h506 : r_q_a <= 20'b01100010000000001000; // 62008 FLAG ---0-,CIN=X_SR
      11'h507 : r_q_a <= 20'b00000000110100001001; // 00D09 LOOP T
      11'h508 : r_q_a <= 20'b11000100001010000000; // C4280 LSHB.
      11'h509 : r_q_a <= 20'b01100001101000001001; // 61A09 FLAG *--0*,CIN=C_FLG
      11'h50A : r_q_a <= 20'b00111110000110011011; // 3E19B JUMP Write_DnB
      11'h50B : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h50C : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h50D : r_q_a <= 20'b00111110010100010000; // 3E510 JUMP ROLB_jmp
      11'h50E : r_q_a <= 20'b10100101000010000000; // A5080 LDB DL[EA1]
      11'h50F : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h510 : r_q_a <= 20'b01100110100000001010; // 6680A FLAG ---00,CIN=N[7]
      11'h511 : r_q_a <= 20'b00000000110100010011; // 00D13 LOOP T
      11'h512 : r_q_a <= 20'b11000100001010000000; // C4280 LSHB.
      11'h513 : r_q_a <= 20'b01100100100000001001; // 64809 FLAG ---0*,CIN=T[7]
      11'h514 : r_q_a <= 20'b00111110000110011011; // 3E19B JUMP Write_DnB
      11'h515 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h516 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h517 : r_q_a <= 20'b00111110010100011010; // 3E51A JUMP ASRW_jmp
      11'h518 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h519 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h51A : r_q_a <= 20'b01100111000000001010; // 6700A FLAG ---00,CIN=N[15]
      11'h51B : r_q_a <= 20'b00000000110100011101; // 00D1D LOOP T
      11'h51C : r_q_a <= 20'b11000100011011000000; // C46C0 RSHW.
      11'h51D : r_q_a <= 20'b01100101001000001001; // 65209 FLAG *--0*,CIN=T[15]
      11'h51E : r_q_a <= 20'b00111110000110011000; // 3E198 JUMP Write_DnW
      11'h51F : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h520 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h521 : r_q_a <= 20'b00111110010100100100; // 3E524 JUMP LSRW_jmp
      11'h522 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h523 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h524 : r_q_a <= 20'b01100000100000001010; // 6080A FLAG ---00,CIN=CLR
      11'h525 : r_q_a <= 20'b00000000110100100111; // 00D27 LOOP T
      11'h526 : r_q_a <= 20'b11000100011011000000; // C46C0 RSHW.
      11'h527 : r_q_a <= 20'b01100000101000001001; // 60A09 FLAG *--0*,CIN=CLR
      11'h528 : r_q_a <= 20'b00111110000110011000; // 3E198 JUMP Write_DnW
      11'h529 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h52A : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h52B : r_q_a <= 20'b00111110010100101110; // 3E52E JUMP ROXRW_jmp
      11'h52C : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h52D : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h52E : r_q_a <= 20'b01100010000000001000; // 62008 FLAG ---0-,CIN=X_SR
      11'h52F : r_q_a <= 20'b00000000110100110001; // 00D31 LOOP T
      11'h530 : r_q_a <= 20'b11000100011011000000; // C46C0 RSHW.
      11'h531 : r_q_a <= 20'b01100001101000001001; // 61A09 FLAG *--0*,CIN=C_FLG
      11'h532 : r_q_a <= 20'b00111110000110011000; // 3E198 JUMP Write_DnW
      11'h533 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h534 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h535 : r_q_a <= 20'b00111110010100111000; // 3E538 JUMP RORW_jmp
      11'h536 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h537 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h538 : r_q_a <= 20'b01100110000000001010; // 6600A FLAG ---00,CIN=N[0]
      11'h539 : r_q_a <= 20'b00000000110100111011; // 00D3B LOOP T
      11'h53A : r_q_a <= 20'b11000100011011000000; // C46C0 RSHW.
      11'h53B : r_q_a <= 20'b01100100000000001001; // 64009 FLAG ---0*,CIN=T[0]
      11'h53C : r_q_a <= 20'b00111110000110011000; // 3E198 JUMP Write_DnW
      11'h53D : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h53E : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h53F : r_q_a <= 20'b00111110010101000010; // 3E542 JUMP ASLW_jmp
      11'h540 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h541 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h542 : r_q_a <= 20'b01100000100000001010; // 6080A FLAG ---00,CIN=CLR
      11'h543 : r_q_a <= 20'b00000000110101000101; // 00D45 LOOP T
      11'h544 : r_q_a <= 20'b11000100011010000000; // C4680 LSHW.
      11'h545 : r_q_a <= 20'b01100000101000000101; // 60A05 FLAG *--**,CIN=CLR
      11'h546 : r_q_a <= 20'b00111110000110011000; // 3E198 JUMP Write_DnW
      11'h547 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h548 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h549 : r_q_a <= 20'b00111110010101001100; // 3E54C JUMP LSLW_jmp
      11'h54A : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h54B : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h54C : r_q_a <= 20'b01100000100000001010; // 6080A FLAG ---00,CIN=CLR
      11'h54D : r_q_a <= 20'b00000000110101001111; // 00D4F LOOP T
      11'h54E : r_q_a <= 20'b11000100011010000000; // C4680 LSHW.
      11'h54F : r_q_a <= 20'b01100000101000001001; // 60A09 FLAG *--0*,CIN=CLR
      11'h550 : r_q_a <= 20'b00111110000110011000; // 3E198 JUMP Write_DnW
      11'h551 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h552 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h553 : r_q_a <= 20'b00111110010101010110; // 3E556 JUMP ROXLW_jmp
      11'h554 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h555 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h556 : r_q_a <= 20'b01100010000000001000; // 62008 FLAG ---0-,CIN=X_SR
      11'h557 : r_q_a <= 20'b00000000110101011001; // 00D59 LOOP T
      11'h558 : r_q_a <= 20'b11000100011010000000; // C4680 LSHW.
      11'h559 : r_q_a <= 20'b01100001101000001001; // 61A09 FLAG *--0*,CIN=C_FLG
      11'h55A : r_q_a <= 20'b00111110000110011000; // 3E198 JUMP Write_DnW
      11'h55B : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h55C : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h55D : r_q_a <= 20'b00111110010101100000; // 3E560 JUMP ROLW_jmp
      11'h55E : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h55F : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h560 : r_q_a <= 20'b01100111000000001010; // 6700A FLAG ---00,CIN=N[15]
      11'h561 : r_q_a <= 20'b00000000110101100011; // 00D63 LOOP T
      11'h562 : r_q_a <= 20'b11000100011010000000; // C4680 LSHW.
      11'h563 : r_q_a <= 20'b01100101000000001001; // 65009 FLAG ---0*,CIN=T[15]
      11'h564 : r_q_a <= 20'b00111110000110011000; // 3E198 JUMP Write_DnW
      11'h565 : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h566 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h567 : r_q_a <= 20'b01100111000000001010; // 6700A FLAG ---00,CIN=N[15]
      11'h568 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h569 : r_q_a <= 20'b00111110010101101110; // 3E56E JUMP ASRL_jmp
      11'h56A : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h56B : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h56C : r_q_a <= 20'b01100111000000001010; // 6700A FLAG ---00,CIN=N[15]
      11'h56D : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h56E : r_q_a <= 20'b00000000110101110000; // 00D70 LOOP T
      11'h56F : r_q_a <= 20'b11000100101011000000; // C4AC0 RSHL.
      11'h570 : r_q_a <= 20'b01100111001000001001; // 67209 FLAG *--0*,CIN=N[15]
      11'h571 : r_q_a <= 20'b00111110000110010011; // 3E193 JUMP Write_DnL
      11'h572 : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h573 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h574 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h575 : r_q_a <= 20'b00111110010101111001; // 3E579 JUMP LSRL_jmp
      11'h576 : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h577 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h578 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h579 : r_q_a <= 20'b01100000100000001010; // 6080A FLAG ---00,CIN=CLR
      11'h57A : r_q_a <= 20'b00000000110101111100; // 00D7C LOOP T
      11'h57B : r_q_a <= 20'b11000100101011000000; // C4AC0 RSHL.
      11'h57C : r_q_a <= 20'b01100000101000001001; // 60A09 FLAG *--0*,CIN=CLR
      11'h57D : r_q_a <= 20'b00111110000110010011; // 3E193 JUMP Write_DnL
      11'h57E : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h57F : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h580 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h581 : r_q_a <= 20'b00111110010110000101; // 3E585 JUMP ROXRL_jmp
      11'h582 : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h583 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h584 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h585 : r_q_a <= 20'b01100010000000001000; // 62008 FLAG ---0-,CIN=X_SR
      11'h586 : r_q_a <= 20'b00000000110110001000; // 00D88 LOOP T
      11'h587 : r_q_a <= 20'b11000100101011000000; // C4AC0 RSHL.
      11'h588 : r_q_a <= 20'b01100001101000001001; // 61A09 FLAG *--0*,CIN=C_FLG
      11'h589 : r_q_a <= 20'b00111110000110010011; // 3E193 JUMP Write_DnL
      11'h58A : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h58B : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h58C : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h58D : r_q_a <= 20'b00111110010110010001; // 3E591 JUMP RORL_jmp
      11'h58E : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h58F : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h590 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h591 : r_q_a <= 20'b01100110000000001010; // 6600A FLAG ---00,CIN=N[0]
      11'h592 : r_q_a <= 20'b00000000110110010100; // 00D94 LOOP T
      11'h593 : r_q_a <= 20'b01100100000000001001; // 64009 FLAG ---0*,CIN=T[0]
      11'h594 : r_q_a <= 20'b11000100101011000000; // C4AC0 RSHL.
      11'h595 : r_q_a <= 20'b00111110000110010011; // 3E193 JUMP Write_DnL
      11'h596 : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h597 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h598 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h599 : r_q_a <= 20'b00111110010110011101; // 3E59D JUMP ASLL_jmp
      11'h59A : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h59B : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h59C : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h59D : r_q_a <= 20'b01100000100000001010; // 6080A FLAG ---00,CIN=CLR
      11'h59E : r_q_a <= 20'b00000000110110100000; // 00DA0 LOOP T
      11'h59F : r_q_a <= 20'b11000100101010000000; // C4A80 LSHL.
      11'h5A0 : r_q_a <= 20'b01100000101000000101; // 60A05 FLAG *--**,CIN=CLR
      11'h5A1 : r_q_a <= 20'b00111110000110010011; // 3E193 JUMP Write_DnL
      11'h5A2 : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h5A3 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h5A4 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h5A5 : r_q_a <= 20'b00111110010110101001; // 3E5A9 JUMP LSLL_jmp
      11'h5A6 : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h5A7 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h5A8 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h5A9 : r_q_a <= 20'b01100000100000001010; // 6080A FLAG ---00,CIN=CLR
      11'h5AA : r_q_a <= 20'b00000000110110101100; // 00DAC LOOP T
      11'h5AB : r_q_a <= 20'b11000100101010000000; // C4A80 LSHL.
      11'h5AC : r_q_a <= 20'b01100000101000001001; // 60A09 FLAG *--0*,CIN=CLR
      11'h5AD : r_q_a <= 20'b00111110000110010011; // 3E193 JUMP Write_DnL
      11'h5AE : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h5AF : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h5B0 : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h5B1 : r_q_a <= 20'b00111110010110110101; // 3E5B5 JUMP ROXLL_jmp
      11'h5B2 : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h5B3 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h5B4 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h5B5 : r_q_a <= 20'b01100010000000001000; // 62008 FLAG ---0-,CIN=X_SR
      11'h5B6 : r_q_a <= 20'b00000000110110111000; // 00DB8 LOOP T
      11'h5B7 : r_q_a <= 20'b11000100101010000000; // C4A80 LSHL.
      11'h5B8 : r_q_a <= 20'b01100001101000001001; // 61A09 FLAG *--0*,CIN=C_FLG
      11'h5B9 : r_q_a <= 20'b00111110000110010011; // 3E193 JUMP Write_DnL
      11'h5BA : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h5BB : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h5BC : r_q_a <= 20'b01100111000000001010; // 6700A FLAG ---00,CIN=N[15]
      11'h5BD : r_q_a <= 20'b10100101010010000100; // A5484 LDW DL[EA2]
      11'h5BE : r_q_a <= 20'b00111110010111000011; // 3E5C3 JUMP ROLL_jmp
      11'h5BF : r_q_a <= 20'b10100101010110000000; // A5580 LDW DH[EA1]
      11'h5C0 : r_q_a <= 20'b10100101010010000000; // A5480 LDW DL[EA1]
      11'h5C1 : r_q_a <= 20'b01100111000000001010; // 6700A FLAG ---00,CIN=N[15]
      11'h5C2 : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h5C3 : r_q_a <= 20'b00000000110111000101; // 00DC5 LOOP T
      11'h5C4 : r_q_a <= 20'b01100111000000001001; // 67009 FLAG ---0*,CIN=N[15]
      11'h5C5 : r_q_a <= 20'b11000100101010000000; // C4A80 LSHL.
      11'h5C6 : r_q_a <= 20'b00111110000110010011; // 3E193 JUMP Write_DnL
      11'h5C7 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h5C8 : r_q_a <= 20'b01100101000000000000; // 65000 FLAG -----,CIN=T[15]
      11'h5C9 : r_q_a <= 20'b11000100011011000000; // C46C0 RSHW.
      11'h5CA : r_q_a <= 20'b01100000101010011001; // 60A99 FLAG ***0*,CIN=CLR
      11'h5CB : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h5CC : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h5CD : r_q_a <= 20'b01100000100000000000; // 60800 FLAG -----,CIN=CLR
      11'h5CE : r_q_a <= 20'b11000100011011000000; // C46C0 RSHW.
      11'h5CF : r_q_a <= 20'b01100000101010011001; // 60A99 FLAG ***0*,CIN=CLR
      11'h5D0 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h5D1 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h5D2 : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h5D3 : r_q_a <= 20'b11000100011011000000; // C46C0 RSHW.
      11'h5D4 : r_q_a <= 20'b01100000101010011001; // 60A99 FLAG ***0*,CIN=CLR
      11'h5D5 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h5D6 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h5D7 : r_q_a <= 20'b01100100000000000000; // 64000 FLAG -----,CIN=T[0]
      11'h5D8 : r_q_a <= 20'b11000100011011000000; // C46C0 RSHW.
      11'h5D9 : r_q_a <= 20'b01100000100010011001; // 60899 FLAG -**0*,CIN=CLR
      11'h5DA : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h5DB : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h5DC : r_q_a <= 20'b01100000100000000000; // 60800 FLAG -----,CIN=CLR
      11'h5DD : r_q_a <= 20'b11000100011010000000; // C4680 LSHW.
      11'h5DE : r_q_a <= 20'b01100000101010010101; // 60A95 FLAG *****,CIN=CLR
      11'h5DF : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h5E0 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h5E1 : r_q_a <= 20'b01100000100000000000; // 60800 FLAG -----,CIN=CLR
      11'h5E2 : r_q_a <= 20'b11000100011010000000; // C4680 LSHW.
      11'h5E3 : r_q_a <= 20'b01100000101010011001; // 60A99 FLAG ***0*,CIN=CLR
      11'h5E4 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h5E5 : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h5E6 : r_q_a <= 20'b01100010000000000000; // 62000 FLAG -----,CIN=X_SR
      11'h5E7 : r_q_a <= 20'b11000100011010000000; // C4680 LSHW.
      11'h5E8 : r_q_a <= 20'b01100000101010011001; // 60A99 FLAG ***0*,CIN=CLR
      11'h5E9 : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h5EA : r_q_a <= 20'b00101110011000000000; // 2E600 CALL EA1_Read_W
      11'h5EB : r_q_a <= 20'b01100101000000000000; // 65000 FLAG -----,CIN=T[15]
      11'h5EC : r_q_a <= 20'b11000100011010000000; // C4680 LSHW.
      11'h5ED : r_q_a <= 20'b01100000100010011001; // 60899 FLAG -**0*,CIN=CLR
      11'h5EE : r_q_a <= 20'b00111110011000110110; // 3E636 JUMP EA1_Update_W
      11'h5EF : r_q_a <= 20'b10000101010010001101; // 8548D LDW EA1J
      11'h5F0 : r_q_a <= 20'b00111111011100110000; // 3F730 JUMP 0730(T)
      11'h5F1 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h5F2 : r_q_a <= 20'b10010101000110000000; // 95180 LDB (EA1); RTS
      11'h5F3 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h5F4 : r_q_a <= 20'b10000101000110000100; // 85184 LDB (EA1)+
      11'h5F5 : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h5F6 : r_q_a <= 20'b00101110011011100010; // 2E6E2 CALL Calc_d16_An_EA1
      11'h5F7 : r_q_a <= 20'b10010101000110000000; // 95180 LDB (EA1); RTS
      11'h5F8 : r_q_a <= 20'b00101110011011101100; // 2E6EC CALL Calc_AbsW_EA1
      11'h5F9 : r_q_a <= 20'b10010101000110000000; // 95180 LDB (EA1); RTS
      11'h5FA : r_q_a <= 20'b00101110011011110001; // 2E6F1 CALL Calc_AbsL_EA1
      11'h5FB : r_q_a <= 20'b10010101000110000000; // 95180 LDB (EA1); RTS
      11'h5FC : r_q_a <= 20'b00101110011011110101; // 2E6F5 CALL Calc_d16_PC_EA1
      11'h5FD : r_q_a <= 20'b10010101000110000000; // 95180 LDB (EA1); RTS
      11'h5FE : r_q_a <= 20'b00101110011011111011; // 2E6FB CALL Calc_d8_PC_Rn_EA1
      11'h5FF : r_q_a <= 20'b10010101000110000000; // 95180 LDB (EA1); RTS
      11'h600 : r_q_a <= 20'b10000101010010001101; // 8548D LDW EA1J
      11'h601 : r_q_a <= 20'b00111111011101000000; // 3F740 JUMP 0740(T)
      11'h602 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h603 : r_q_a <= 20'b10010101010110000000; // 95580 LDW (EA1); RTS
      11'h604 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h605 : r_q_a <= 20'b10000101010110000100; // 85584 LDW (EA1)+
      11'h606 : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h607 : r_q_a <= 20'b00101110011011100010; // 2E6E2 CALL Calc_d16_An_EA1
      11'h608 : r_q_a <= 20'b10010101010110000000; // 95580 LDW (EA1); RTS
      11'h609 : r_q_a <= 20'b00101110011011101100; // 2E6EC CALL Calc_AbsW_EA1
      11'h60A : r_q_a <= 20'b10010101010110000000; // 95580 LDW (EA1); RTS
      11'h60B : r_q_a <= 20'b00101110011011110001; // 2E6F1 CALL Calc_AbsL_EA1
      11'h60C : r_q_a <= 20'b10010101010110000000; // 95580 LDW (EA1); RTS
      11'h60D : r_q_a <= 20'b00101110011011110101; // 2E6F5 CALL Calc_d16_PC_EA1
      11'h60E : r_q_a <= 20'b10010101010110000000; // 95580 LDW (EA1); RTS
      11'h60F : r_q_a <= 20'b00101110011011111011; // 2E6FB CALL Calc_d8_PC_Rn_EA1
      11'h610 : r_q_a <= 20'b10010101010110000000; // 95580 LDW (EA1); RTS
      11'h611 : r_q_a <= 20'b10000101010010001101; // 8548D LDW EA1J
      11'h612 : r_q_a <= 20'b00111111011101010000; // 3F750 JUMP 0750(T)
      11'h613 : r_q_a <= 20'b10100101010110000010; // A5582 LDW RH[EA1]
      11'h614 : r_q_a <= 20'b10110101010010000010; // B5482 LDW RL[EA1]; RTS
      11'h615 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h616 : r_q_a <= 20'b00111110011101011110; // 3E75E JUMP EA1_RL
      11'h617 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h618 : r_q_a <= 20'b10000101010110000100; // 85584 LDW (EA1)+
      11'h619 : r_q_a <= 20'b10000101010110000100; // 85584 LDW (EA1)+
      11'h61A : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h61B : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h61C : r_q_a <= 20'b10000101010110001000; // 85588 LDW -(EA1)
      11'h61D : r_q_a <= 20'b10000101010110001000; // 85588 LDW -(EA1)
      11'h61E : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h61F : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h620 : r_q_a <= 20'b00101110011011100010; // 2E6E2 CALL Calc_d16_An_EA1
      11'h621 : r_q_a <= 20'b00111110011101011110; // 3E75E JUMP EA1_RL
      11'h622 : r_q_a <= 20'b00101110011011101100; // 2E6EC CALL Calc_AbsW_EA1
      11'h623 : r_q_a <= 20'b00111110011101011110; // 3E75E JUMP EA1_RL
      11'h624 : r_q_a <= 20'b00101110011011110001; // 2E6F1 CALL Calc_AbsL_EA1
      11'h625 : r_q_a <= 20'b00111110011101011110; // 3E75E JUMP EA1_RL
      11'h626 : r_q_a <= 20'b00101110011011110101; // 2E6F5 CALL Calc_d16_PC_EA1
      11'h627 : r_q_a <= 20'b00111110011101011110; // 3E75E JUMP EA1_RL
      11'h628 : r_q_a <= 20'b00101110011011111011; // 2E6FB CALL Calc_d8_PC_Rn_EA1
      11'h629 : r_q_a <= 20'b00111110011101011110; // 3E75E JUMP EA1_RL
      11'h62A : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h62B : r_q_a <= 20'b10100011010101001100; // A354C STW TMP1H
      11'h62C : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h62D : r_q_a <= 20'b10100011010001001100; // A344C STW TMP1L
      11'h62E : r_q_a <= 20'b00101110011000010001; // 2E611 CALL EA1_Read_L
      11'h62F : r_q_a <= 20'b10110101010010001100; // B548C LDW TMP1L; RTS
      11'h630 : r_q_a <= 20'b10000101010010001101; // 8548D LDW EA1J
      11'h631 : r_q_a <= 20'b00111111011101100000; // 3F760 JUMP 0760(T)
      11'h632 : r_q_a <= 20'b00110110011101110000; // 36770 JUMP EA7,EA1_WB_Reg
      11'h633 : r_q_a <= 20'b00110101011000110101; // 35635 JUMP EA4,EA1_UpdB_An
      11'h634 : r_q_a <= 20'b10010011000101000001; // 93141 STB (EA2); RTS
      11'h635 : r_q_a <= 20'b10010011000101000100; // 93144 STB (EA1)+; RTS
      11'h636 : r_q_a <= 20'b00110110011110000000; // 36780 JUMP EA7,EA1_WW_Reg
      11'h637 : r_q_a <= 20'b00110101011000111001; // 35639 JUMP EA4,EA1_UpdW_An
      11'h638 : r_q_a <= 20'b10010011010101000001; // 93541 STW (EA2); RTS
      11'h639 : r_q_a <= 20'b10010011010101000000; // 93540 STW (EA1); RTS
      11'h63A : r_q_a <= 20'b00110110011001010001; // 36651 JUMP EA7,EA1_WL_Reg
      11'h63B : r_q_a <= 20'b00110101011110011010; // 3579A JUMP EA4,EA1_WL
      11'h63C : r_q_a <= 20'b00111110011111001010; // 3E7CA JUMP EA2_WL
      11'h63D : r_q_a <= 20'b10000101010010001101; // 8548D LDW EA1J
      11'h63E : r_q_a <= 20'b00111111011101110000; // 3F770 JUMP 0770(T)
      11'h63F : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h640 : r_q_a <= 20'b10010011000101000000; // 93140 STB (EA1); RTS
      11'h641 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h642 : r_q_a <= 20'b10000011000101000100; // 83144 STB (EA1)+
      11'h643 : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h644 : r_q_a <= 20'b00101110011011100010; // 2E6E2 CALL Calc_d16_An_EA1
      11'h645 : r_q_a <= 20'b10010011000101000000; // 93140 STB (EA1); RTS
      11'h646 : r_q_a <= 20'b10000101010010001101; // 8548D LDW EA1J
      11'h647 : r_q_a <= 20'b00111111011110000000; // 3F780 JUMP 0780(T)
      11'h648 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h649 : r_q_a <= 20'b10010011010101000000; // 93540 STW (EA1); RTS
      11'h64A : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h64B : r_q_a <= 20'b10000011010101000100; // 83544 STW (EA1)+
      11'h64C : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h64D : r_q_a <= 20'b00101110011011100010; // 2E6E2 CALL Calc_d16_An_EA1
      11'h64E : r_q_a <= 20'b10010011010101000000; // 93540 STW (EA1); RTS
      11'h64F : r_q_a <= 20'b10000101010010001101; // 8548D LDW EA1J
      11'h650 : r_q_a <= 20'b00111111011110010000; // 3F790 JUMP 0790(T)
      11'h651 : r_q_a <= 20'b10100011010101000010; // A3542 STW RH[EA1]
      11'h652 : r_q_a <= 20'b10110011010001000010; // B3442 STW RL[EA1]; RTS
      11'h653 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h654 : r_q_a <= 20'b00111110011110011010; // 3E79A JUMP EA1_WL
      11'h655 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h656 : r_q_a <= 20'b10000011010101000100; // 83544 STW (EA1)+
      11'h657 : r_q_a <= 20'b10000011010101000100; // 83544 STW (EA1)+
      11'h658 : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h659 : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h65A : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h65B : r_q_a <= 20'b10000011010101001000; // 83548 STW -(EA1)
      11'h65C : r_q_a <= 20'b10000011010101001000; // 83548 STW -(EA1)
      11'h65D : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h65E : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h65F : r_q_a <= 20'b10000101000110000101; // 85185 LDB (EA2)+
      11'h660 : r_q_a <= 20'b00111110011100001010; // 3E70A JUMP Set_An_EA2
      11'h661 : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h662 : r_q_a <= 20'b10000101000110001001; // 85189 LDB -(EA2)
      11'h663 : r_q_a <= 20'b00111110011100001010; // 3E70A JUMP Set_An_EA2
      11'h664 : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h665 : r_q_a <= 20'b10000101010110000101; // 85585 LDW (EA2)+
      11'h666 : r_q_a <= 20'b00111110011100001010; // 3E70A JUMP Set_An_EA2
      11'h667 : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h668 : r_q_a <= 20'b10000101010110001001; // 85589 LDW -(EA2)
      11'h669 : r_q_a <= 20'b00111110011100001010; // 3E70A JUMP Set_An_EA2
      11'h66A : r_q_a <= 20'b10000101010010001110; // 8548E LDW EA2J
      11'h66B : r_q_a <= 20'b00111111011110100000; // 3F7A0 JUMP 07A0(T)
      11'h66C : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h66D : r_q_a <= 20'b10010011000101000001; // 93141 STB (EA2); RTS
      11'h66E : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h66F : r_q_a <= 20'b10000011000101000101; // 83145 STB (EA2)+
      11'h670 : r_q_a <= 20'b00111110011100001010; // 3E70A JUMP Set_An_EA2
      11'h671 : r_q_a <= 20'b00101110011100010111; // 2E717 CALL Calc_d16_An_EA2
      11'h672 : r_q_a <= 20'b10010011000101000001; // 93141 STB (EA2); RTS
      11'h673 : r_q_a <= 20'b10000101010010001110; // 8548E LDW EA2J
      11'h674 : r_q_a <= 20'b00111111011110110000; // 3F7B0 JUMP 07B0(T)
      11'h675 : r_q_a <= 20'b01100101000000000000; // 65000 FLAG -----,CIN=T[15]
      11'h676 : r_q_a <= 20'b10100011010001000101; // A3445 STW AL[EA2]
      11'h677 : r_q_a <= 20'b11000101010000110001; // C5431 EXTW
      11'h678 : r_q_a <= 20'b10110011010101000101; // B3545 STW AH[EA2]; RTS
      11'h679 : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h67A : r_q_a <= 20'b10010011010101000001; // 93541 STW (EA2); RTS
      11'h67B : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h67C : r_q_a <= 20'b10000011010101000101; // 83545 STW (EA2)+
      11'h67D : r_q_a <= 20'b00111110011100001010; // 3E70A JUMP Set_An_EA2
      11'h67E : r_q_a <= 20'b00101110011100010111; // 2E717 CALL Calc_d16_An_EA2
      11'h67F : r_q_a <= 20'b10010011010101000001; // 93541 STW (EA2); RTS
      11'h680 : r_q_a <= 20'b10000101010010001110; // 8548E LDW EA2J
      11'h681 : r_q_a <= 20'b00111111011111000000; // 3F7C0 JUMP 07C0(T)
      11'h682 : r_q_a <= 20'b10100011010101000110; // A3546 STW RH[EA2]
      11'h683 : r_q_a <= 20'b10110011010001000110; // B3446 STW RL[EA2]; RTS
      11'h684 : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h685 : r_q_a <= 20'b00111110011111001010; // 3E7CA JUMP EA2_WL
      11'h686 : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h687 : r_q_a <= 20'b10000011010101000101; // 83545 STW (EA2)+
      11'h688 : r_q_a <= 20'b10000011010101000101; // 83545 STW (EA2)+
      11'h689 : r_q_a <= 20'b00111110011100001010; // 3E70A JUMP Set_An_EA2
      11'h68A : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h68B : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h68C : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h68D : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h68E : r_q_a <= 20'b00111110011100001010; // 3E70A JUMP Set_An_EA2
      11'h68F : r_q_a <= 20'b10000101010010001000; // 85488 LDW IMM
      11'h690 : r_q_a <= 20'b01100101000000000000; // 65000 FLAG -----,CIN=T[15]
      11'h691 : r_q_a <= 20'b11000011011000001010; // C360A ADDW.
      11'h692 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h693 : r_q_a <= 20'b11000101010000110001; // C5431 EXTW
      11'h694 : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h695 : r_q_a <= 20'b11010011100000011010; // D381A ADDCL; RTS
      11'h696 : r_q_a <= 20'b10100101010010001010; // A548A LDW RL[EXT]
      11'h697 : r_q_a <= 20'b01100101000000000000; // 65000 FLAG -----,CIN=T[15]
      11'h698 : r_q_a <= 20'b11000011011000001010; // C360A ADDW.
      11'h699 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h69A : r_q_a <= 20'b00110111011010011110; // 3769E JUMP EXT11,LongRn
      11'h69B : r_q_a <= 20'b11000101010000110001; // C5431 EXTW
      11'h69C : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h69D : r_q_a <= 20'b11010011100000011010; // D381A ADDCL; RTS
      11'h69E : r_q_a <= 20'b10100101010110001010; // A558A LDW RH[EXT]
      11'h69F : r_q_a <= 20'b01100001000000000000; // 61000 FLAG -----,CIN=C_ADD
      11'h6A0 : r_q_a <= 20'b11010011100000011010; // D381A ADDCL; RTS
      11'h6A1 : r_q_a <= 20'b00101110011010110010; // 2E6B2 CALL SP_to_EA2
      11'h6A2 : r_q_a <= 20'b10000101010010000100; // 85484 LDW PCL
      11'h6A3 : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h6A4 : r_q_a <= 20'b10000101010010000101; // 85485 LDW PCH
      11'h6A5 : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h6A6 : r_q_a <= 20'b10000101010010001111; // 8548F LDW SR
      11'h6A7 : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h6A8 : r_q_a <= 20'b00111110011010101110; // 3E6AE JUMP EA2_to_SP
      11'h6A9 : r_q_a <= 20'b00101110011010110010; // 2E6B2 CALL SP_to_EA2
      11'h6AA : r_q_a <= 20'b10000101010010000100; // 85484 LDW PCL
      11'h6AB : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h6AC : r_q_a <= 20'b10000101010010000101; // 85485 LDW PCH
      11'h6AD : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h6AE : r_q_a <= 20'b10000101010010000011; // 85483 LDW EA2H
      11'h6AF : r_q_a <= 20'b10100011010101000011; // A3543 STW A7H
      11'h6B0 : r_q_a <= 20'b10000101010010000010; // 85482 LDW EA2L
      11'h6B1 : r_q_a <= 20'b10110011010001000011; // B3443 STW A7L; RTS
      11'h6B2 : r_q_a <= 20'b10100101010110000011; // A5583 LDW A7H
      11'h6B3 : r_q_a <= 20'b10000011010001000011; // 83443 STW EA2H
      11'h6B4 : r_q_a <= 20'b10100101010010000011; // A5483 LDW A7L
      11'h6B5 : r_q_a <= 20'b10010011010001000010; // 93442 STW EA2L; RTS
      11'h6B6 : r_q_a <= 20'b10100101010110000011; // A5583 LDW A7H
      11'h6B7 : r_q_a <= 20'b10100011010101001110; // A354E STW USPH
      11'h6B8 : r_q_a <= 20'b10100101010010000011; // A5483 LDW A7L
      11'h6B9 : r_q_a <= 20'b10110011010001001110; // B344E STW USPL; RTS
      11'h6BA : r_q_a <= 20'b10100101010110000011; // A5583 LDW A7H
      11'h6BB : r_q_a <= 20'b10100011010101001111; // A354F STW SSPH
      11'h6BC : r_q_a <= 20'b10100101010010000011; // A5483 LDW A7L
      11'h6BD : r_q_a <= 20'b10110011010001001111; // B344F STW SSPL; RTS
      11'h6BE : r_q_a <= 20'b00111100011010111010; // 3C6BA JUMP S_SR,A7_to_SSP
      11'h6BF : r_q_a <= 20'b00101110011010110110; // 2E6B6 CALL A7_to_USP
      11'h6C0 : r_q_a <= 20'b10100101010110001111; // A558F LDW SSPH
      11'h6C1 : r_q_a <= 20'b10100011010101000011; // A3543 STW A7H
      11'h6C2 : r_q_a <= 20'b10100101010010001111; // A548F LDW SSPL
      11'h6C3 : r_q_a <= 20'b10110011010001000011; // B3443 STW A7L; RTS
      11'h6C4 : r_q_a <= 20'b10100101010110001110; // A558E LDW USPH
      11'h6C5 : r_q_a <= 20'b10100011010101000011; // A3543 STW A7H
      11'h6C6 : r_q_a <= 20'b10100101010010001110; // A548E LDW USPL
      11'h6C7 : r_q_a <= 20'b10110011010001000011; // B3443 STW A7L; RTS
      11'h6C8 : r_q_a <= 20'b00101110011010111010; // 2E6BA CALL A7_to_SSP
      11'h6C9 : r_q_a <= 20'b00111100111011000100; // 3CEC4 JUMPN S_SR,USP_to_A7
      11'h6CA : r_q_a <= 20'b11010000010001011000; // D0458 NOP; RTS
      11'h6CB : r_q_a <= 20'b10000101010010001111; // 8548F LDW SR
      11'h6CC : r_q_a <= 20'b01000111111111111111; // 47FFF LIT #7FFF
      11'h6CD : r_q_a <= 20'b11000011010001001010; // C344A ANDW
      11'h6CE : r_q_a <= 20'b01000010000000000000; // 42000 LIT #2000
      11'h6CF : r_q_a <= 20'b11010011010001011010; // D345A ORW; RTS
      11'h6D0 : r_q_a <= 20'b10000011010001001111; // 8344F STW SR
      11'h6D1 : r_q_a <= 20'b10000101010110000111; // 85587 LDW (VEC)+
      11'h6D2 : r_q_a <= 20'b10000011010001000101; // 83445 STW PCH
      11'h6D3 : r_q_a <= 20'b10000101010110000111; // 85587 LDW (VEC)+
      11'h6D4 : r_q_a <= 20'b10000011010001000100; // 83444 STW PCL
      11'h6D5 : r_q_a <= 20'b01000000000001100000; // 40060 LIT #0060
      11'h6D6 : r_q_a <= 20'b10010011010001000110; // 93446 STW VECL; RTS
      11'h6D7 : r_q_a <= 20'b10100101010110000001; // A5581 LDW AH[EA1]
      11'h6D8 : r_q_a <= 20'b10100101010010000001; // A5481 LDW AL[EA1]
      11'h6D9 : r_q_a <= 20'b00111110011010001111; // 3E68F JUMP AddOffs
      11'h6DA : r_q_a <= 20'b10100101010010000001; // A5481 LDW AL[EA1]
      11'h6DB : r_q_a <= 20'b10000011010001000000; // 83440 STW EA1L
      11'h6DC : r_q_a <= 20'b10100101010110000001; // A5581 LDW AH[EA1]
      11'h6DD : r_q_a <= 20'b10010011010001000001; // 93441 STW EA1H; RTS
      11'h6DE : r_q_a <= 20'b10000101010010000000; // 85480 LDW EA1L
      11'h6DF : r_q_a <= 20'b10100011010001000001; // A3441 STW AL[EA1]
      11'h6E0 : r_q_a <= 20'b10000101010010000001; // 85481 LDW EA1H
      11'h6E1 : r_q_a <= 20'b10110011010101000001; // B3541 STW AH[EA1]; RTS
      11'h6E2 : r_q_a <= 20'b10000000010110001010; // 8058A FTW (PC)+
      11'h6E3 : r_q_a <= 20'b00101110011011010111; // 2E6D7 CALL Add_Offs_An_EA1
      11'h6E4 : r_q_a <= 20'b10000011010001000001; // 83441 STW EA1H
      11'h6E5 : r_q_a <= 20'b10010011010001000000; // 93440 STW EA1L; RTS
      11'h6E6 : r_q_a <= 20'b10000000010110000110; // 80586 FTE (PC)+
      11'h6E7 : r_q_a <= 20'b00101110011011010111; // 2E6D7 CALL Add_Offs_An_EA1
      11'h6E8 : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h6E9 : r_q_a <= 20'b00101110011010010110; // 2E696 CALL Add_Ext_Rn
      11'h6EA : r_q_a <= 20'b10000011010001000001; // 83441 STW EA1H
      11'h6EB : r_q_a <= 20'b10010011010001000000; // 93440 STW EA1L; RTS
      11'h6EC : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h6ED : r_q_a <= 20'b01100101000000000000; // 65000 FLAG -----,CIN=T[15]
      11'h6EE : r_q_a <= 20'b11000101010000110001; // C5431 EXTW
      11'h6EF : r_q_a <= 20'b10000011010001000001; // 83441 STW EA1H
      11'h6F0 : r_q_a <= 20'b10010011010001000000; // 93440 STW EA1L; RTS
      11'h6F1 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h6F2 : r_q_a <= 20'b10000011010001000001; // 83441 STW EA1H
      11'h6F3 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h6F4 : r_q_a <= 20'b10010011010001000000; // 93440 STW EA1L; RTS
      11'h6F5 : r_q_a <= 20'b10000101010010000101; // 85485 LDW PCH
      11'h6F6 : r_q_a <= 20'b10000101010010000100; // 85484 LDW PCL
      11'h6F7 : r_q_a <= 20'b10000000010110001010; // 8058A FTW (PC)+
      11'h6F8 : r_q_a <= 20'b00101110011010001111; // 2E68F CALL AddOffs
      11'h6F9 : r_q_a <= 20'b10000011010001000001; // 83441 STW EA1H
      11'h6FA : r_q_a <= 20'b10010011010001000000; // 93440 STW EA1L; RTS
      11'h6FB : r_q_a <= 20'b10000101010010000101; // 85485 LDW PCH
      11'h6FC : r_q_a <= 20'b10000101010010000100; // 85484 LDW PCL
      11'h6FD : r_q_a <= 20'b10000000010110000110; // 80586 FTE (PC)+
      11'h6FE : r_q_a <= 20'b00101110011010001111; // 2E68F CALL AddOffs
      11'h6FF : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h700 : r_q_a <= 20'b00101110011010010110; // 2E696 CALL Add_Ext_Rn
      11'h701 : r_q_a <= 20'b10000011010001000001; // 83441 STW EA1H
      11'h702 : r_q_a <= 20'b10010011010001000000; // 93440 STW EA1L; RTS
      11'h703 : r_q_a <= 20'b10100101010110000101; // A5585 LDW AH[EA2]
      11'h704 : r_q_a <= 20'b10100101010010000101; // A5485 LDW AL[EA2]
      11'h705 : r_q_a <= 20'b00111110011010001111; // 3E68F JUMP AddOffs
      11'h706 : r_q_a <= 20'b10100101010010000101; // A5485 LDW AL[EA2]
      11'h707 : r_q_a <= 20'b10000011010001000010; // 83442 STW EA2L
      11'h708 : r_q_a <= 20'b10100101010110000101; // A5585 LDW AH[EA2]
      11'h709 : r_q_a <= 20'b10010011010001000011; // 93443 STW EA2H; RTS
      11'h70A : r_q_a <= 20'b10000101010010000010; // 85482 LDW EA2L
      11'h70B : r_q_a <= 20'b10100011010001000101; // A3445 STW AL[EA2]
      11'h70C : r_q_a <= 20'b10000101010010000011; // 85483 LDW EA2H
      11'h70D : r_q_a <= 20'b10110011010101000101; // B3545 STW AH[EA2]; RTS
      11'h70E : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h70F : r_q_a <= 20'b01100101000000000000; // 65000 FLAG -----,CIN=T[15]
      11'h710 : r_q_a <= 20'b11000101010000110001; // C5431 EXTW
      11'h711 : r_q_a <= 20'b10000011010001000011; // 83443 STW EA2H
      11'h712 : r_q_a <= 20'b10010011010001000010; // 93442 STW EA2L; RTS
      11'h713 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h714 : r_q_a <= 20'b10000011010001000011; // 83443 STW EA2H
      11'h715 : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h716 : r_q_a <= 20'b10010011010001000010; // 93442 STW EA2L; RTS
      11'h717 : r_q_a <= 20'b10000000010110001010; // 8058A FTW (PC)+
      11'h718 : r_q_a <= 20'b00101110011100000011; // 2E703 CALL Add_Offs_An_EA2
      11'h719 : r_q_a <= 20'b10000011010001000011; // 83443 STW EA2H
      11'h71A : r_q_a <= 20'b10010011010001000010; // 93442 STW EA2L; RTS
      11'h71B : r_q_a <= 20'b10000000010110000110; // 80586 FTE (PC)+
      11'h71C : r_q_a <= 20'b00101110011100000011; // 2E703 CALL Add_Offs_An_EA2
      11'h71D : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h71E : r_q_a <= 20'b00101110011010010110; // 2E696 CALL Add_Ext_Rn
      11'h71F : r_q_a <= 20'b10000011010001000011; // 83443 STW EA2H
      11'h720 : r_q_a <= 20'b10010011010001000010; // 93442 STW EA2L; RTS
      11'h721 : r_q_a <= 20'b10000101010010000101; // 85485 LDW PCH
      11'h722 : r_q_a <= 20'b10000101010010000100; // 85484 LDW PCL
      11'h723 : r_q_a <= 20'b10000000010110001010; // 8058A FTW (PC)+
      11'h724 : r_q_a <= 20'b00101110011010001111; // 2E68F CALL AddOffs
      11'h725 : r_q_a <= 20'b10000011010001000011; // 83443 STW EA2H
      11'h726 : r_q_a <= 20'b10010011010001000010; // 93442 STW EA2L; RTS
      11'h727 : r_q_a <= 20'b10000101010010000101; // 85485 LDW PCH
      11'h728 : r_q_a <= 20'b10000101010010000100; // 85484 LDW PCL
      11'h729 : r_q_a <= 20'b10000000010110000110; // 80586 FTE (PC)+
      11'h72A : r_q_a <= 20'b00101110011010001111; // 2E68F CALL AddOffs
      11'h72B : r_q_a <= 20'b11000100010001010010; // C4452 SWAP
      11'h72C : r_q_a <= 20'b00101110011010010110; // 2E696 CALL Add_Ext_Rn
      11'h72D : r_q_a <= 20'b10000011010001000011; // 83443 STW EA2H
      11'h72E : r_q_a <= 20'b10010011010001000010; // 93442 STW EA2L; RTS
      11'h72F : r_q_a <= 20'b00000000000000000000; // 00000 
      11'h730 : r_q_a <= 20'b10110101000010000010; // B5082 LDB RL[EA1]; RTS
      11'h731 : r_q_a <= 20'b00111110000000000000; // 3E000 JUMP 0000
      11'h732 : r_q_a <= 20'b00111110010111110001; // 3E5F1 JUMP EA1_RB_An
      11'h733 : r_q_a <= 20'b00111110010111110011; // 3E5F3 JUMP EA1_RB_An_Inc
      11'h734 : r_q_a <= 20'b00111110011100111101; // 3E73D JUMP EA1_RB_An_Dec
      11'h735 : r_q_a <= 20'b00111110010111110110; // 3E5F6 JUMP EA1_RB_d16_An
      11'h736 : r_q_a <= 20'b00101110011011100110; // 2E6E6 CALL Calc_d8_An_Rn_EA1
      11'h737 : r_q_a <= 20'b10010101000110000000; // 95180 LDB (EA1); RTS
      11'h738 : r_q_a <= 20'b00111110010111111000; // 3E5F8 JUMP EA1_RB_AbsW
      11'h739 : r_q_a <= 20'b00111110010111111010; // 3E5FA JUMP EA1_RB_AbsL
      11'h73A : r_q_a <= 20'b00111110010111111100; // 3E5FC JUMP EA1_RB_d16_PC
      11'h73B : r_q_a <= 20'b00111110010111111110; // 3E5FE JUMP EA1_RB_d8_PC_Rn
      11'h73C : r_q_a <= 20'b10010101010110001010; // 9558A LDW (PC)+; RTS
      11'h73D : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h73E : r_q_a <= 20'b10000101000110001000; // 85188 LDB -(EA1)
      11'h73F : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h740 : r_q_a <= 20'b10110101010010000010; // B5482 LDW RL[EA1]; RTS
      11'h741 : r_q_a <= 20'b10110101010010000010; // B5482 LDW RL[EA1]; RTS
      11'h742 : r_q_a <= 20'b00111110011000000010; // 3E602 JUMP EA1_RW_An
      11'h743 : r_q_a <= 20'b00111110011000000100; // 3E604 JUMP EA1_RW_An_Inc
      11'h744 : r_q_a <= 20'b00111110011101001101; // 3E74D JUMP EA1_RW_An_Dec
      11'h745 : r_q_a <= 20'b00111110011000000111; // 3E607 JUMP EA1_RW_d16_An
      11'h746 : r_q_a <= 20'b00101110011011100110; // 2E6E6 CALL Calc_d8_An_Rn_EA1
      11'h747 : r_q_a <= 20'b10010101010110000000; // 95580 LDW (EA1); RTS
      11'h748 : r_q_a <= 20'b00111110011000001001; // 3E609 JUMP EA1_RW_AbsW
      11'h749 : r_q_a <= 20'b00111110011000001011; // 3E60B JUMP EA1_RW_AbsL
      11'h74A : r_q_a <= 20'b00111110011000001101; // 3E60D JUMP EA1_RW_d16_PC
      11'h74B : r_q_a <= 20'b00111110011000001111; // 3E60F JUMP EA1_RW_d8_PC_Rn
      11'h74C : r_q_a <= 20'b10010101010110001010; // 9558A LDW (PC)+; RTS
      11'h74D : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h74E : r_q_a <= 20'b10000101010110001000; // 85588 LDW -(EA1)
      11'h74F : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h750 : r_q_a <= 20'b00111110011000010011; // 3E613 JUMP EA1_RL_Reg
      11'h751 : r_q_a <= 20'b00111110011000010011; // 3E613 JUMP EA1_RL_Reg
      11'h752 : r_q_a <= 20'b00111110011000010101; // 3E615 JUMP EA1_RL_An
      11'h753 : r_q_a <= 20'b00111110011000010111; // 3E617 JUMP EA1_RL_An_Inc
      11'h754 : r_q_a <= 20'b00111110011000011011; // 3E61B JUMP EA1_RL_An_Dec
      11'h755 : r_q_a <= 20'b00111110011000100000; // 3E620 JUMP EA1_RL_d16_An
      11'h756 : r_q_a <= 20'b00101110011011100110; // 2E6E6 CALL Calc_d8_An_Rn_EA1
      11'h757 : r_q_a <= 20'b00111110011101011110; // 3E75E JUMP EA1_RL
      11'h758 : r_q_a <= 20'b00111110011000100010; // 3E622 JUMP EA1_RL_AbsW
      11'h759 : r_q_a <= 20'b00111110011000100100; // 3E624 JUMP EA1_RL_AbsL
      11'h75A : r_q_a <= 20'b00111110011000100110; // 3E626 JUMP EA1_RL_d16_PC
      11'h75B : r_q_a <= 20'b00111110011000101000; // 3E628 JUMP EA1_RL_d8_PC_Rn
      11'h75C : r_q_a <= 20'b10000101010110001010; // 8558A LDW (PC)+
      11'h75D : r_q_a <= 20'b10010101010110001010; // 9558A LDW (PC)+; RTS
      11'h75E : r_q_a <= 20'b10000101010110000100; // 85584 LDW (EA1)+
      11'h75F : r_q_a <= 20'b10010101010110000000; // 95580 LDW (EA1); RTS
      11'h760 : r_q_a <= 20'b00111110000000000000; // 3E000 JUMP 0000
      11'h761 : r_q_a <= 20'b00111110000000000000; // 3E000 JUMP 0000
      11'h762 : r_q_a <= 20'b00111110011011011010; // 3E6DA JUMP Get_An_EA1
      11'h763 : r_q_a <= 20'b00111110011011011010; // 3E6DA JUMP Get_An_EA1
      11'h764 : r_q_a <= 20'b00111110011011011010; // 3E6DA JUMP Get_An_EA1
      11'h765 : r_q_a <= 20'b00111110011011100010; // 3E6E2 JUMP Calc_d16_An_EA1
      11'h766 : r_q_a <= 20'b00111110011011100110; // 3E6E6 JUMP Calc_d8_An_Rn_EA1
      11'h767 : r_q_a <= 20'b00111110000000000000; // 3E000 JUMP 0000
      11'h768 : r_q_a <= 20'b00111110011011101100; // 3E6EC JUMP Calc_AbsW_EA1
      11'h769 : r_q_a <= 20'b00111110011011110001; // 3E6F1 JUMP Calc_AbsL_EA1
      11'h76A : r_q_a <= 20'b00111110011011110101; // 3E6F5 JUMP Calc_d16_PC_EA1
      11'h76B : r_q_a <= 20'b00111110011011111011; // 3E6FB JUMP Calc_d8_PC_Rn_EA1
      11'h76C : r_q_a <= 20'b00111110000000000000; // 3E000 JUMP 0000
      11'h76D : r_q_a <= 20'b00111110000000000000; // 3E000 JUMP 0000
      11'h76E : r_q_a <= 20'b00111110000000000000; // 3E000 JUMP 0000
      11'h76F : r_q_a <= 20'b00111110000000000000; // 3E000 JUMP 0000
      11'h770 : r_q_a <= 20'b10110011000001000010; // B3042 STB RL[EA1]; RTS
      11'h771 : r_q_a <= 20'b00111110000000000000; // 3E000 JUMP 0000
      11'h772 : r_q_a <= 20'b00111110011000111111; // 3E63F JUMP EA1_WB_An
      11'h773 : r_q_a <= 20'b00111110011001000001; // 3E641 JUMP EA1_WB_An_Inc
      11'h774 : r_q_a <= 20'b00111110011101111101; // 3E77D JUMP EA1_WB_An_Dec
      11'h775 : r_q_a <= 20'b00111110011001000100; // 3E644 JUMP EA1_WB_d16_An
      11'h776 : r_q_a <= 20'b00101110011011100110; // 2E6E6 CALL Calc_d8_An_Rn_EA1
      11'h777 : r_q_a <= 20'b10010011000101000000; // 93140 STB (EA1); RTS
      11'h778 : r_q_a <= 20'b00111110011101111011; // 3E77B JUMP EA1_WB_AbsW
      11'h779 : r_q_a <= 20'b00101110011011110001; // 2E6F1 CALL Calc_AbsL_EA1
      11'h77A : r_q_a <= 20'b10010011000101000000; // 93140 STB (EA1); RTS
      11'h77B : r_q_a <= 20'b00101110011011101100; // 2E6EC CALL Calc_AbsW_EA1
      11'h77C : r_q_a <= 20'b10010011000101000000; // 93140 STB (EA1); RTS
      11'h77D : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h77E : r_q_a <= 20'b10000011000101001000; // 83148 STB -(EA1)
      11'h77F : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h780 : r_q_a <= 20'b10110011010001000010; // B3442 STW RL[EA1]; RTS
      11'h781 : r_q_a <= 20'b00111110000000000000; // 3E000 JUMP 0000
      11'h782 : r_q_a <= 20'b00111110011001001000; // 3E648 JUMP EA1_WW_An
      11'h783 : r_q_a <= 20'b00111110011001001010; // 3E64A JUMP EA1_WW_An_Inc
      11'h784 : r_q_a <= 20'b00111110011110001101; // 3E78D JUMP EA1_WW_An_Dec
      11'h785 : r_q_a <= 20'b00111110011001001101; // 3E64D JUMP EA1_WW_d16_An
      11'h786 : r_q_a <= 20'b00101110011011100110; // 2E6E6 CALL Calc_d8_An_Rn_EA1
      11'h787 : r_q_a <= 20'b10010011010101000000; // 93540 STW (EA1); RTS
      11'h788 : r_q_a <= 20'b00111110011110001011; // 3E78B JUMP EA1_WW_AbsW
      11'h789 : r_q_a <= 20'b00101110011011110001; // 2E6F1 CALL Calc_AbsL_EA1
      11'h78A : r_q_a <= 20'b10010011010101000000; // 93540 STW (EA1); RTS
      11'h78B : r_q_a <= 20'b00101110011011101100; // 2E6EC CALL Calc_AbsW_EA1
      11'h78C : r_q_a <= 20'b10010011010101000000; // 93540 STW (EA1); RTS
      11'h78D : r_q_a <= 20'b00101110011011011010; // 2E6DA CALL Get_An_EA1
      11'h78E : r_q_a <= 20'b10000011010101001000; // 83548 STW -(EA1)
      11'h78F : r_q_a <= 20'b00111110011011011110; // 3E6DE JUMP Set_An_EA1
      11'h790 : r_q_a <= 20'b00111110011001010001; // 3E651 JUMP EA1_WL_Reg
      11'h791 : r_q_a <= 20'b00111110011001010001; // 3E651 JUMP EA1_WL_Reg
      11'h792 : r_q_a <= 20'b00111110011001010011; // 3E653 JUMP EA1_WL_An
      11'h793 : r_q_a <= 20'b00111110011001010101; // 3E655 JUMP EA1_WL_An_Inc
      11'h794 : r_q_a <= 20'b00111110011001011001; // 3E659 JUMP EA1_WL_An_Dec
      11'h795 : r_q_a <= 20'b00111110011110011100; // 3E79C JUMP EA1_WL_d16_An
      11'h796 : r_q_a <= 20'b00101110011011100110; // 2E6E6 CALL Calc_d8_An_Rn_EA1
      11'h797 : r_q_a <= 20'b00111110011110011010; // 3E79A JUMP EA1_WL
      11'h798 : r_q_a <= 20'b00111110011110011110; // 3E79E JUMP EA1_WL_AbsW
      11'h799 : r_q_a <= 20'b00101110011011110001; // 2E6F1 CALL Calc_AbsL_EA1
      11'h79A : r_q_a <= 20'b10000011010101000100; // 83544 STW (EA1)+
      11'h79B : r_q_a <= 20'b10010011010101000000; // 93540 STW (EA1); RTS
      11'h79C : r_q_a <= 20'b00101110011011100010; // 2E6E2 CALL Calc_d16_An_EA1
      11'h79D : r_q_a <= 20'b00111110011110011010; // 3E79A JUMP EA1_WL
      11'h79E : r_q_a <= 20'b00101110011011101100; // 2E6EC CALL Calc_AbsW_EA1
      11'h79F : r_q_a <= 20'b00111110011110011010; // 3E79A JUMP EA1_WL
      11'h7A0 : r_q_a <= 20'b10110011000001000100; // B3044 STB DL[EA2]; RTS
      11'h7A1 : r_q_a <= 20'b00111110000000000000; // 3E000 JUMP 0000
      11'h7A2 : r_q_a <= 20'b00111110011001101100; // 3E66C JUMP EA2_WB_An
      11'h7A3 : r_q_a <= 20'b00111110011001101110; // 3E66E JUMP EA2_WB_An_Inc
      11'h7A4 : r_q_a <= 20'b00111110011110101101; // 3E7AD JUMP EA2_WB_An_Dec
      11'h7A5 : r_q_a <= 20'b00111110011001110001; // 3E671 JUMP EA2_WB_d16_An
      11'h7A6 : r_q_a <= 20'b00101110011100011011; // 2E71B CALL Calc_d8_An_Rn_EA2
      11'h7A7 : r_q_a <= 20'b10010011000101000001; // 93141 STB (EA2); RTS
      11'h7A8 : r_q_a <= 20'b00111110011110101011; // 3E7AB JUMP EA2_WB_AbsW
      11'h7A9 : r_q_a <= 20'b00101110011100010011; // 2E713 CALL Calc_AbsL_EA2
      11'h7AA : r_q_a <= 20'b10010011000101000001; // 93141 STB (EA2); RTS
      11'h7AB : r_q_a <= 20'b00101110011100001110; // 2E70E CALL Calc_AbsW_EA2
      11'h7AC : r_q_a <= 20'b10010011000101000001; // 93141 STB (EA2); RTS
      11'h7AD : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h7AE : r_q_a <= 20'b10000011000101001001; // 83149 STB -(EA2)
      11'h7AF : r_q_a <= 20'b00111110011100001010; // 3E70A JUMP Set_An_EA2
      11'h7B0 : r_q_a <= 20'b10110011010001000110; // B3446 STW RL[EA2]; RTS
      11'h7B1 : r_q_a <= 20'b00111110011001110101; // 3E675 JUMP EA2_WW_AReg
      11'h7B2 : r_q_a <= 20'b00111110011001111001; // 3E679 JUMP EA2_WW_An
      11'h7B3 : r_q_a <= 20'b00111110011001111011; // 3E67B JUMP EA2_WW_An_Inc
      11'h7B4 : r_q_a <= 20'b00111110011110111101; // 3E7BD JUMP EA2_WW_An_Dec
      11'h7B5 : r_q_a <= 20'b00111110011001111110; // 3E67E JUMP EA2_WW_d16_An
      11'h7B6 : r_q_a <= 20'b00101110011100011011; // 2E71B CALL Calc_d8_An_Rn_EA2
      11'h7B7 : r_q_a <= 20'b10010011010101000001; // 93541 STW (EA2); RTS
      11'h7B8 : r_q_a <= 20'b00111110011110111011; // 3E7BB JUMP EA2_WW_AbsW
      11'h7B9 : r_q_a <= 20'b00101110011100010011; // 2E713 CALL Calc_AbsL_EA2
      11'h7BA : r_q_a <= 20'b10010011010101000001; // 93541 STW (EA2); RTS
      11'h7BB : r_q_a <= 20'b00101110011100001110; // 2E70E CALL Calc_AbsW_EA2
      11'h7BC : r_q_a <= 20'b10010011010101000001; // 93541 STW (EA2); RTS
      11'h7BD : r_q_a <= 20'b00101110011100000110; // 2E706 CALL Get_An_EA2
      11'h7BE : r_q_a <= 20'b10000011010101001001; // 83549 STW -(EA2)
      11'h7BF : r_q_a <= 20'b00111110011100001010; // 3E70A JUMP Set_An_EA2
      11'h7C0 : r_q_a <= 20'b00111110011010000010; // 3E682 JUMP EA2_WL_Reg
      11'h7C1 : r_q_a <= 20'b00111110011010000010; // 3E682 JUMP EA2_WL_Reg
      11'h7C2 : r_q_a <= 20'b00111110011010000100; // 3E684 JUMP EA2_WL_An
      11'h7C3 : r_q_a <= 20'b00111110011010000110; // 3E686 JUMP EA2_WL_An_Inc
      11'h7C4 : r_q_a <= 20'b00111110011010001010; // 3E68A JUMP EA2_WL_An_Dec
      11'h7C5 : r_q_a <= 20'b00111110011111001100; // 3E7CC JUMP EA2_WL_d16_An
      11'h7C6 : r_q_a <= 20'b00101110011100011011; // 2E71B CALL Calc_d8_An_Rn_EA2
      11'h7C7 : r_q_a <= 20'b00111110011111001010; // 3E7CA JUMP EA2_WL
      11'h7C8 : r_q_a <= 20'b00111110011111001110; // 3E7CE JUMP EA2_WL_AbsW
      11'h7C9 : r_q_a <= 20'b00101110011100010011; // 2E713 CALL Calc_AbsL_EA2
      11'h7CA : r_q_a <= 20'b10000011010101000101; // 83545 STW (EA2)+
      11'h7CB : r_q_a <= 20'b10010011010101000001; // 93541 STW (EA2); RTS
      11'h7CC : r_q_a <= 20'b00101110011100010111; // 2E717 CALL Calc_d16_An_EA2
      11'h7CD : r_q_a <= 20'b00111110011111001010; // 3E7CA JUMP EA2_WL
      11'h7CE : r_q_a <= 20'b00101110011100001110; // 2E70E CALL Calc_AbsW_EA2
      11'h7CF : r_q_a <= 20'b00111110011111001010; // 3E7CA JUMP EA2_WL
      11'h7D0 : r_q_a <= 20'b11000000010001011000; // C0458 NOP
      11'h7D1 : r_q_a <= 20'b11000000010001011000; // C0458 NOP
      11'h7D2 : r_q_a <= 20'b11000000010001011000; // C0458 NOP
      11'h7D3 : r_q_a <= 20'b11000000010001011000; // C0458 NOP
      11'h7D4 : r_q_a <= 20'b11000000010001011000; // C0458 NOP
      11'h7D5 : r_q_a <= 20'b11000000010001011000; // C0458 NOP
      11'h7D6 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7D7 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7D8 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7D9 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7DA : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7DB : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7DC : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7DD : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7DE : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7DF : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7E0 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7E1 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7E2 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7E3 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7E4 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7E5 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7E6 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7E7 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7E8 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7E9 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7EA : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7EB : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7EC : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7ED : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7EE : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7EF : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7F0 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7F1 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7F2 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7F3 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7F4 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7F5 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7F6 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7F7 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7F8 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7F9 : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7FA : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7FB : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7FC : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7FD : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7FE : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
      11'h7FF : r_q_a <= 20'b01000000000000000000; // 40000 LIT #0000
    endcase
  end
end

assign q_a = r_q_a;

// Port B (read/write)
always@(posedge clock) begin
  r_q_b <= r_mem_blk[address_b][15:0];
  if (wren_b[0]) r_mem_blk[address_b][7:0]  <= data_b[7:0];
  if (wren_b[1]) r_mem_blk[address_b][15:8] <= data_b[15:8];
end

assign q_b = r_q_b;

endmodule
