module decode_rom
(
  input         clock,
  input   [7:0] address,
  output [35:0] q
);

reg  [35:0] r_q;

always@(posedge clock) begin
  case(address)
    8'h00 : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h01 : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h02 : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h03 : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h04 : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h05 : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h06 : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h07 : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h08 : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h09 : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h0A : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h0B : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h0C : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h0D : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h0E : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h0F : r_q <= 36'b001000000010_000000_000000_1110_00000000; // 202, +0, +0
    8'h10 : r_q <= 36'b001000000100_000000_000000_1110_00000000; // 204, +0, +0
    8'h11 : r_q <= 36'b001000000100_000000_000000_1110_00000000; // 204, +0, +0
    8'h12 : r_q <= 36'b001000000100_000000_000000_1110_00000000; // 204, +0, +0
    8'h13 : r_q <= 36'b001000000100_000000_000000_1110_00000000; // 204, +0, +0
    8'h14 : r_q <= 36'b001000000100_000000_000000_1110_00000000; // 204, +0, +0
    8'h15 : r_q <= 36'b001000000100_000000_000000_1110_00000000; // 204, +0, +0
    8'h16 : r_q <= 36'b001000000100_000000_000000_1110_00000000; // 204, +0, +0
    8'h17 : r_q <= 36'b001000000100_000000_000000_1110_00000000; // 204, +0, +0
    8'h18 : r_q <= 36'b001000010001_000000_000000_1110_00000000; // 211, +0, +0
    8'h19 : r_q <= 36'b001000010001_000000_000000_1110_00000000; // 211, +0, +0
    8'h1A : r_q <= 36'b001000010001_000000_000000_1110_00000000; // 211, +0, +0
    8'h1B : r_q <= 36'b001000010001_000000_000000_1110_00000000; // 211, +0, +0
    8'h1C : r_q <= 36'b001000010001_000000_000000_1110_00000000; // 211, +0, +0
    8'h1D : r_q <= 36'b001000010001_000000_000000_1110_00000000; // 211, +0, +0
    8'h1E : r_q <= 36'b001000010001_000000_000000_1110_00000000; // 211, +0, +0
    8'h1F : r_q <= 36'b001000010001_000000_000000_1110_00000000; // 211, +0, +0
    8'h20 : r_q <= 36'b001000011101_000000_000000_1110_00000000; // 21D, +0, +0
    8'h21 : r_q <= 36'b001000011101_000000_000000_1110_00000000; // 21D, +0, +0
    8'h22 : r_q <= 36'b001000011101_000000_000000_1110_00000000; // 21D, +0, +0
    8'h23 : r_q <= 36'b001000011101_000000_000000_1110_00000000; // 21D, +0, +0
    8'h24 : r_q <= 36'b001000011101_000000_000000_1110_00000000; // 21D, +0, +0
    8'h25 : r_q <= 36'b001000011101_000000_000000_1110_00000000; // 21D, +0, +0
    8'h26 : r_q <= 36'b001000011101_000000_000000_1110_00000000; // 21D, +0, +0
    8'h27 : r_q <= 36'b001000011101_000000_000000_1110_00000000; // 21D, +0, +0
    8'h28 : r_q <= 36'b001000100001_000000_000000_1110_00000000; // 221, +0, +0
    8'h29 : r_q <= 36'b001000100001_000000_000000_1110_00000000; // 221, +0, +0
    8'h2A : r_q <= 36'b001000100001_000000_000000_1110_00000000; // 221, +0, +0
    8'h2B : r_q <= 36'b001000100001_000000_000000_1110_00000000; // 221, +0, +0
    8'h2C : r_q <= 36'b001000100001_000000_000000_1110_00000000; // 221, +0, +0
    8'h2D : r_q <= 36'b001000100001_000000_000000_1110_00000000; // 221, +0, +0
    8'h2E : r_q <= 36'b001000100001_000000_000000_1110_00000000; // 221, +0, +0
    8'h2F : r_q <= 36'b001000100001_000000_000000_1110_00000000; // 221, +0, +0
    8'h30 : r_q <= 36'b000000000000_000000_000000_1110_00000000; // 000, +0, +0
    8'h31 : r_q <= 36'b001000000001_000000_000000_1110_00000000; // 201, +0, +0
    8'h32 : r_q <= 36'b001000100101_000000_000000_1110_00000000; // 225, +0, +0
    8'h33 : r_q <= 36'b001000101001_000000_000000_1110_00000000; // 229, +0, +0
    8'h34 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h35 : r_q <= 36'b001000101110_000000_000000_1110_00000000; // 22E, +0, +0
    8'h36 : r_q <= 36'b001000110100_000000_000000_1110_00000000; // 234, +0, +0
    8'h37 : r_q <= 36'b001000110111_000000_000000_1110_00000000; // 237, +0, +0
    8'h38 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h39 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h3A : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h3B : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h3C : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h3D : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h3E : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h3F : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h40 : r_q <= 36'b000001000110_000000_000101_1011_00000000; // 046, +0, +5
    8'h41 : r_q <= 36'b000001001111_000000_000101_1011_00000000; // 04F, +0, +5
    8'h42 : r_q <= 36'b000001011001_000000_000000_0011_00000000; // 059, +0, +0
    8'h43 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h44 : r_q <= 36'b000001100000_000000_000101_1011_00000000; // 060, +0, +5
    8'h45 : r_q <= 36'b000001101001_000000_000101_1011_00000000; // 069, +0, +5
    8'h46 : r_q <= 36'b000001110011_000000_000000_0011_00000000; // 073, +0, +0
    8'h47 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h48 : r_q <= 36'b000001111010_000000_000000_0011_00000000; // 07A, +0, +0
    8'h49 : r_q <= 36'b000001111111_000000_000000_0011_00000000; // 07F, +0, +0
    8'h4A : r_q <= 36'b000010000100_000000_000000_0011_00000000; // 084, +0, +0
    8'h4B : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h4C : r_q <= 36'b000010001100_000000_000000_0011_00000000; // 08C, +0, +0
    8'h4D : r_q <= 36'b000010010001_000000_000000_0011_00000000; // 091, +0, +0
    8'h4E : r_q <= 36'b000010010110_000000_000000_0011_00000000; // 096, +0, +0
    8'h4F : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h50 : r_q <= 36'b000010011110_001011_001011_1010_00000000; // 09E, +11, +11
    8'h51 : r_q <= 36'b000010110010_000100_000100_0011_00000000; // 0B2, +4, +4
    8'h52 : r_q <= 36'b000010111111_000100_000100_0011_00000000; // 0BF, +4, +4
    8'h53 : r_q <= 36'b000011001100_000100_000100_0011_00000000; // 0CC, +4, +4
    8'h54 : r_q <= 36'b000011011001_000000_000101_1011_00000000; // 0D9, +0, +5
    8'h55 : r_q <= 36'b000011100010_000000_000101_1011_00000000; // 0E2, +0, +5
    8'h56 : r_q <= 36'b000011101100_000000_000000_0011_00000000; // 0EC, +0, +0
    8'h57 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h58 : r_q <= 36'b000011110011_000000_000000_0011_00000000; // 0F3, +0, +0
    8'h59 : r_q <= 36'b000011111000_000000_000000_0011_00000000; // 0F8, +0, +0
    8'h5A : r_q <= 36'b000011111101_000000_000000_0011_00000000; // 0FD, +0, +0
    8'h5B : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h5C : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h5D : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h5E : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h5F : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h60 : r_q <= 36'b000101000100_000000_000000_0011_00000000; // 144, +0, +0
    8'h61 : r_q <= 36'b000101001001_000000_000000_0011_00000000; // 149, +0, +0
    8'h62 : r_q <= 36'b000101001110_000000_000000_0011_00000000; // 14E, +0, +0
    8'h63 : r_q <= 36'b000101010110_000000_000000_0011_00000000; // 156, +0, +0
    8'h64 : r_q <= 36'b000101011000_000000_000000_0011_00000000; // 158, +0, +0
    8'h65 : r_q <= 36'b000101011011_000000_000000_0011_00000000; // 15B, +0, +0
    8'h66 : r_q <= 36'b000101011110_000000_000000_0011_00000000; // 15E, +0, +0
    8'h67 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h68 : r_q <= 36'b000101100010_000000_000000_0011_00000000; // 162, +0, +0
    8'h69 : r_q <= 36'b000101100110_000000_000000_0011_00000000; // 166, +0, +0
    8'h6A : r_q <= 36'b000101101010_000000_000000_0011_00000000; // 16A, +0, +0
    8'h6B : r_q <= 36'b000101110001_000000_000000_1100_00000000; // 171, +0, +0
    8'h6C : r_q <= 36'b000101110011_000000_000000_0011_00000000; // 173, +0, +0
    8'h6D : r_q <= 36'b000101110111_000000_000000_0011_00000000; // 177, +0, +0
    8'h6E : r_q <= 36'b000101111011_000000_000000_0011_00000000; // 17B, +0, +0
    8'h6F : r_q <= 36'b000110000001_000000_000000_1100_00000000; // 181, +0, +0
    8'h70 : r_q <= 36'b000110000100_000000_000000_0011_00000000; // 184, +0, +0
    8'h71 : r_q <= 36'b000110001001_000111_000000_1000_00000000; // 189, +7, +0
    8'h72 : r_q <= 36'b000110011110_010001_001000_0001_00000000; // 19E, +17, +8
    8'h73 : r_q <= 36'b000110111000_010101_001010_0001_00000000; // 1B8, +21, +10
    8'h74 : r_q <= 36'b000111010011_000000_000000_0011_00000000; // 1D3, +0, +0
    8'h75 : r_q <= 36'b000111010111_000000_000000_0011_00000000; // 1D7, +0, +0
    8'h76 : r_q <= 36'b000111011011_000000_000000_0011_00000000; // 1DB, +0, +0
    8'h77 : r_q <= 36'b000111100001_000000_000000_0011_00000000; // 1E1, +0, +0
    8'h78 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h79 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h7A : r_q <= 36'b000111100111_000000_001100_1001_00000000; // 1E7, +0, +12
    8'h7B : r_q <= 36'b000111110101_000000_001010_1001_00000000; // 1F5, +0, +10
    8'h7C : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h7D : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'h7E : r_q <= 36'b001000111011_000000_000000_0111_00000000; // 23B, +0, +0
    8'h7F : r_q <= 36'b001001000001_000000_000000_0111_00000000; // 241, +0, +0
    8'h80 : r_q <= 36'b010011001000_000000_000000_1110_00000000; // 4C8, +0, +0
    8'h81 : r_q <= 36'b010011010010_000000_000000_1110_00000000; // 4D2, +0, +0
    8'h82 : r_q <= 36'b010011011100_000000_000000_1110_00000000; // 4DC, +0, +0
    8'h83 : r_q <= 36'b010011100110_000000_000000_1110_00000000; // 4E6, +0, +0
    8'h84 : r_q <= 36'b010011000101_000000_000000_1110_00000000; // 4C5, +0, +0
    8'h85 : r_q <= 36'b010011001111_000000_000000_1110_00000000; // 4CF, +0, +0
    8'h86 : r_q <= 36'b010011011001_000000_000000_1110_00000000; // 4D9, +0, +0
    8'h87 : r_q <= 36'b010011100011_000000_000000_1110_00000000; // 4E3, +0, +0
    8'h88 : r_q <= 36'b010011110000_000000_000000_1110_00000000; // 4F0, +0, +0
    8'h89 : r_q <= 36'b010011111010_000000_000000_1110_00000000; // 4FA, +0, +0
    8'h8A : r_q <= 36'b010100000100_000000_000000_1110_00000000; // 504, +0, +0
    8'h8B : r_q <= 36'b010100001110_000000_000000_1110_00000000; // 50E, +0, +0
    8'h8C : r_q <= 36'b010011101101_000000_000000_1110_00000000; // 4ED, +0, +0
    8'h8D : r_q <= 36'b010011110111_000000_000000_1110_00000000; // 4F7, +0, +0
    8'h8E : r_q <= 36'b010100000001_000000_000000_1110_00000000; // 501, +0, +0
    8'h8F : r_q <= 36'b010100001011_000000_000000_1110_00000000; // 50B, +0, +0
    8'h90 : r_q <= 36'b010100011000_000000_000000_1110_00000000; // 518, +0, +0
    8'h91 : r_q <= 36'b010100100010_000000_000000_1110_00000000; // 522, +0, +0
    8'h92 : r_q <= 36'b010100101100_000000_000000_1110_00000000; // 52C, +0, +0
    8'h93 : r_q <= 36'b010100110110_000000_000000_1110_00000000; // 536, +0, +0
    8'h94 : r_q <= 36'b010100010101_000000_000000_1110_00000000; // 515, +0, +0
    8'h95 : r_q <= 36'b010100011111_000000_000000_1110_00000000; // 51F, +0, +0
    8'h96 : r_q <= 36'b010100101001_000000_000000_1110_00000000; // 529, +0, +0
    8'h97 : r_q <= 36'b010100110011_000000_000000_1110_00000000; // 533, +0, +0
    8'h98 : r_q <= 36'b010101000000_000000_000000_1110_00000000; // 540, +0, +0
    8'h99 : r_q <= 36'b010101001010_000000_000000_1110_00000000; // 54A, +0, +0
    8'h9A : r_q <= 36'b010101010100_000000_000000_1110_00000000; // 554, +0, +0
    8'h9B : r_q <= 36'b010101011110_000000_000000_1110_00000000; // 55E, +0, +0
    8'h9C : r_q <= 36'b010100111101_000000_000000_1110_00000000; // 53D, +0, +0
    8'h9D : r_q <= 36'b010101000111_000000_000000_1110_00000000; // 547, +0, +0
    8'h9E : r_q <= 36'b010101010001_000000_000000_1110_00000000; // 551, +0, +0
    8'h9F : r_q <= 36'b010101011011_000000_000000_1110_00000000; // 55B, +0, +0
    8'hA0 : r_q <= 36'b010101101010_000000_000000_1110_00000000; // 56A, +0, +0
    8'hA1 : r_q <= 36'b010101110110_000000_000000_1110_00000000; // 576, +0, +0
    8'hA2 : r_q <= 36'b010110000010_000000_000000_1110_00000000; // 582, +0, +0
    8'hA3 : r_q <= 36'b010110001110_000000_000000_1110_00000000; // 58E, +0, +0
    8'hA4 : r_q <= 36'b010101100101_000000_000000_1110_00000000; // 565, +0, +0
    8'hA5 : r_q <= 36'b010101110010_000000_000000_1110_00000000; // 572, +0, +0
    8'hA6 : r_q <= 36'b010101111110_000000_000000_1110_00000000; // 57E, +0, +0
    8'hA7 : r_q <= 36'b010110001010_000000_000000_1110_00000000; // 58A, +0, +0
    8'hA8 : r_q <= 36'b010110011010_000000_000000_1110_00000000; // 59A, +0, +0
    8'hA9 : r_q <= 36'b010110100110_000000_000000_1110_00000000; // 5A6, +0, +0
    8'hAA : r_q <= 36'b010110110010_000000_000000_1110_00000000; // 5B2, +0, +0
    8'hAB : r_q <= 36'b010110111111_000000_000000_1110_00000000; // 5BF, +0, +0
    8'hAC : r_q <= 36'b010110010110_000000_000000_1110_00000000; // 596, +0, +0
    8'hAD : r_q <= 36'b010110100010_000000_000000_1110_00000000; // 5A2, +0, +0
    8'hAE : r_q <= 36'b010110101110_000000_000000_1110_00000000; // 5AE, +0, +0
    8'hAF : r_q <= 36'b010110111010_000000_000000_1110_00000000; // 5BA, +0, +0
    8'hB0 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'hB1 : r_q <= 36'b000100110001_000000_000000_1100_00000000; // 131, +0, +0
    8'hB2 : r_q <= 36'b000100110101_000110_000000_1101_00000000; // 135, +6, +0
    8'hB3 : r_q <= 36'b000100111110_000100_000000_1101_00000000; // 13E, +4, +0
    8'hB4 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'hB5 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'hB6 : r_q <= 36'b001010100100_000111_000000_1110_00000000; // 2A4, +7, +0
    8'hB7 : r_q <= 36'b001010110101_000000_000000_1110_00000000; // 2B5, +0, +0
    8'hB8 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'hB9 : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'hBA : r_q <= 36'b000000110100_000000_000000_1110_00000000; // 034, +0, +0
    8'hBB : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'hBC : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'hBD : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'hBE : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'hBF : r_q <= 36'b000000110010_000000_000000_1110_00000000; // 032, +0, +0
    8'hC0 : r_q <= 36'b001010111011_000000_000000_1100_00000000; // 2BB, +0, +0
    8'hC1 : r_q <= 36'b001011100101_000000_000000_1100_00000000; // 2E5, +0, +0
    8'hC2 : r_q <= 36'b001011101101_000000_000000_1100_00000000; // 2ED, +0, +0
    8'hC3 : r_q <= 36'b001011111000_000000_000000_1100_00000000; // 2F8, +0, +0
    8'hC4 : r_q <= 36'b001010111101_000110_001011_0101_00000000; // 2BD, +6, +11
    8'hC5 : r_q <= 36'b001011100111_000000_000000_0010_00000000; // 2E7, +0, +0
    8'hC6 : r_q <= 36'b001011101111_000000_000000_0010_00000000; // 2EF, +0, +0
    8'hC7 : r_q <= 36'b001100010100_000000_000000_1100_00000000; // 314, +0, +0
    8'hC8 : r_q <= 36'b001100110111_000000_000000_1100_00000000; // 337, +0, +0
    8'hC9 : r_q <= 36'b001101001101_000000_000000_1101_00000000; // 34D, +0, +0
    8'hCA : r_q <= 36'b001101100011_000000_000000_1101_00000000; // 363, +0, +0
    8'hCB : r_q <= 36'b001110001111_000000_000000_1101_00000000; // 38F, +0, +0
    8'hCC : r_q <= 36'b001100111100_000101_001011_0101_00000000; // 33C, +5, +11
    8'hCD : r_q <= 36'b001101010010_000101_001011_0101_00000000; // 352, +5, +11
    8'hCE : r_q <= 36'b001101101100_001001_010100_0101_00000000; // 36C, +9, +20
    8'hCF : r_q <= 36'b001110011010_000000_000000_1101_00000000; // 39A, +0, +0
    8'hD0 : r_q <= 36'b001001010111_000000_000000_0011_00000000; // 257, +0, +0
    8'hD1 : r_q <= 36'b001001011100_000000_010000_0101_00000000; // 25C, +0, +16
    8'hD2 : r_q <= 36'b001001100001_000000_001011_0101_00000000; // 261, +0, +11
    8'hD3 : r_q <= 36'b001010010011_000000_000101_0101_00000000; // 293, +0, +5
    8'hD4 : r_q <= 36'b001001110101_000000_000000_0011_00000000; // 275, +0, +0
    8'hD5 : r_q <= 36'b001001111010_000000_010000_0101_00000000; // 27A, +0, +16
    8'hD6 : r_q <= 36'b001001111111_000000_001011_0101_00000000; // 27F, +0, +11
    8'hD7 : r_q <= 36'b001010010011_000000_000101_0101_00000000; // 293, +0, +5
    8'hD8 : r_q <= 36'b001110011100_000000_000000_1100_00000000; // 39C, +0, +0
    8'hD9 : r_q <= 36'b001110100001_000000_000000_1101_00000000; // 3A1, +0, +0
    8'hDA : r_q <= 36'b001110100110_000000_000000_1101_00000000; // 3A6, +0, +0
    8'hDB : r_q <= 36'b001110101111_000000_000000_1101_00000000; // 3AF, +0, +0
    8'hDC : r_q <= 36'b001110111011_000000_000101_0101_00000000; // 3BB, +0, +5
    8'hDD : r_q <= 36'b001111000101_000000_000101_0101_00000000; // 3C5, +0, +5
    8'hDE : r_q <= 36'b001111001111_000000_001000_0101_00000000; // 3CF, +0, +8
    8'hDF : r_q <= 36'b001111100101_000000_000000_1101_00000000; // 3E5, +0, +0
    8'hE0 : r_q <= 36'b001111100111_000000_000000_1100_00000000; // 3E7, +0, +0
    8'hE1 : r_q <= 36'b010000011000_000000_000000_1100_00000000; // 418, +0, +0
    8'hE2 : r_q <= 36'b010000110000_000000_000000_1100_00000000; // 430, +0, +0
    8'hE3 : r_q <= 36'b010001000011_000000_000000_1100_00000000; // 443, +0, +0
    8'hE4 : r_q <= 36'b001111101001_000110_001011_0101_00000000; // 3E9, +6, +11
    8'hE5 : r_q <= 36'b010000011010_000110_001110_0101_00000000; // 41A, +6, +14
    8'hE6 : r_q <= 36'b010000110010_000000_001001_0100_00000000; // 432, +0, +9
    8'hE7 : r_q <= 36'b010001010111_000000_000000_1100_00000000; // 457, +0, +0
    8'hE8 : r_q <= 36'b010001101010_000000_000000_1100_00000000; // 46A, +0, +0
    8'hE9 : r_q <= 36'b010001111110_000000_000000_1101_00000000; // 47E, +0, +0
    8'hEA : r_q <= 36'b010010010010_000000_000000_1101_00000000; // 492, +0, +0
    8'hEB : r_q <= 36'b010010111000_000000_000000_1101_00000000; // 4B8, +0, +0
    8'hEC : r_q <= 36'b010001101100_000110_001100_0101_00000000; // 46C, +6, +12
    8'hED : r_q <= 36'b010010000000_000110_001100_0101_00000000; // 480, +6, +12
    8'hEE : r_q <= 36'b010010010100_001010_010101_0101_00000000; // 494, +10, +21
    8'hEF : r_q <= 36'b010011000011_000000_000000_1101_00000000; // 4C3, +0, +0
    8'hF0 : r_q <= 36'b010111000111_000000_000000_0010_00000000; // 5C7, +0, +0
    8'hF1 : r_q <= 36'b010111011011_000000_000000_0010_00000000; // 5DB, +0, +0
    8'hF2 : r_q <= 36'b010111001100_000000_000000_0010_00000000; // 5CC, +0, +0
    8'hF3 : r_q <= 36'b010111100000_000000_000000_0010_00000000; // 5E0, +0, +0
    8'hF4 : r_q <= 36'b010111010001_000000_000000_0010_00000000; // 5D1, +0, +0
    8'hF5 : r_q <= 36'b010111100101_000000_000000_0010_00000000; // 5E5, +0, +0
    8'hF6 : r_q <= 36'b010111010110_000000_000000_0010_00000000; // 5D6, +0, +0
    8'hF7 : r_q <= 36'b010111101010_000000_000000_0010_00000000; // 5EA, +0, +0
    8'hF8 : r_q <= 36'b000100000101_000010_000100_1101_00000000; // 105, +2, +4
    8'hF9 : r_q <= 36'b000100001011_000010_000110_0101_00000000; // 10B, +2, +6
    8'hFA : r_q <= 36'b000100011010_000010_000110_0101_00000000; // 11A, +2, +6
    8'hFB : r_q <= 36'b000100100010_000010_000110_0101_00000000; // 122, +2, +6
    8'hFC : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'hFD : r_q <= 36'b000000111010_000000_000000_0000_00000000; // 03A, +0, +0
    8'hFE : r_q <= 36'b001001000011_000000_000000_1100_00000000; // 243, +0, +0
    8'hFF : r_q <= 36'b001001010010_000000_000000_0111_00000000; // 252, +0, +0
  endcase
end

endmodule
